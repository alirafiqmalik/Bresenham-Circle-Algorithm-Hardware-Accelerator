module vga_demo(CLOCK_50, SW, KEY_N,
				VGA_R, VGA_G, VGA_B,
				VGA_HS, VGA_VS, VGA_BLANK, VGA_SYNC, VGA_CLK,
				HEX0_N,HEX1_N);
	
	input CLOCK_50;	
	input [9:0] SW;
	input [3:0] KEY_N;
	output [7:0] VGA_R;
	output [7:0] VGA_G;
	output [7:0] VGA_B;
	output VGA_HS;
	output VGA_VS;
	
	output VGA_BLANK;
	output VGA_SYNC;
	output VGA_CLK;	


output [6:0]HEX0_N,HEX1_N;


	

	wire [7:0] x;
	wire [6:0] y;
	

	
	wire [7:0] vga_x;
   wire [6:0] vga_y;
	wire [2:0]vga_colour;	
	wire vga_plot;
	
  //  Bresenham_circle T3T (CLOCK_50,KEY_N,SW,x,y,vga_x,vga_y,vga_plot,vga_colour);	
	// Bresenham_circle  (CLOCK_50,KEY_N,SW,lockingkeyinput,vga_colour,vga_plot,vga_x,vga_y)
  Bresenham_circle Bresenham_circle_init (CLOCK_50,KEY_N,SW,lockingkeyinput,vga_colour,vga_plot,vga_x,vga_y);	

  wire [127:0] lockingkeyinput;
	// assign lockingkeyinput=128'b10101010111110001110011111101001000001001010000100010100011111010111100001001000101110011111101100101000111000010111111001100011;
	wire [3:0] address;
	hexto7segment H0(address,HEX0_N);
	hexto7segment H1({3'b0,address[3]},HEX1_N);

memory_with_timer my_memory (
    .clk(CLOCK_50),
    .reset(1'b1),
    .count_up_key(KEY_N[1]),
    .count_down_key(KEY_N[2]),
    .address(address),
    .data_out(lockingkeyinput)
);

	

	vga_adapter VGA(
			.resetn(KEY_N[3]),
			.clock(CLOCK_50),
			.colour(vga_colour),
			.x(vga_x),
			.y(vga_y),
			.plot(vga_plot),
			/* Signals for the DAC to drive the monitor. */
			.VGA_R(VGA_R),
			.VGA_G(VGA_G),
			.VGA_B(VGA_B),
			.VGA_HS(VGA_HS),
			.VGA_VS(VGA_VS),
			.VGA_BLANK(VGA_BLANK),
			.VGA_SYNC(VGA_SYNC),
			.VGA_CLK(VGA_CLK));
		defparam VGA.RESOLUTION = "160x120";//"320x240";
		defparam VGA.MONOCHROME = "FALSE";
		defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
		defparam VGA.BACKGROUND_IMAGE = "image.colour.mif";
		defparam VGA.USING_DE1 = "TRUE";
		
endmodule
	


module hexto7segment(input [3:0]x,output reg [6:0]z);
	always @(x)
	case (x)
		4'h0 : z = 7'b1000000;
		4'h1 : z = 7'b1111001;
		4'h2 : z = 7'b0100100;
		4'h3 : z = 7'b0110000;
		4'h4 : z = 7'b0011001;
		4'h5 : z = 7'b0010010;
		4'h6 : z = 7'b0000010;
		4'h7 : z = 7'b1111000;
		4'h8 : z = 7'b0000000;
		4'h9 : z = 7'b0010000;
		4'hA : z = 7'b0001000;
		4'hB : z = 7'b0000011;
		4'hC : z = 7'b1000110;
		4'hD : z = 7'b0100001;
		4'hE : z = 7'b0000110;
		4'hF : z = 7'b0001110;
		
	default:z= 7'b1111111; 
	endcase
endmodule



module memory_with_timer (
    clk,
    reset,
    count_up_key,
    count_down_key,
    address,
    data_out);

    parameter n = 4; // Number of address bits
    parameter m = 128; // Number of memory bits per address
    

    input clk;
    input reset;
    input count_up_key;
    input count_down_key;
    output [n-1:0] address;
    output [m-1:0] data_out;

    reg [n-1:0] address_reg;
    reg [m-1:0] memory [0:2**n-1];

		reg [25:0] count;

    // Initialize memory with initial values
    initial 
      begin
			// integer i;
      $readmemb("keys.txt", memory);//Reading and assiging initial values to RAM from "instruction1.txt" file
        // for (i = 0; i < (2**n); i=i+1) begin
        //     memory[i] = i % (2**m);
        // end
    end

    // Assign outputs
    assign address = address_reg;
    assign data_out = memory[address_reg];

    // Count-up and count-down logic
    always @ (posedge clk,negedge reset) begin
        if (!reset) begin
            address_reg = 5;
						count=0;
        end else if(count==26'd25000000) begin
						count=0;
            if (!count_up_key & count_down_key) begin
                address_reg = address_reg + 1;
            end 
						else if (!count_down_key & count_up_key) begin
                address_reg = address_reg - 1;
            end
        end
				else count=count+1;
    end

endmodule

// 128'b10101010111110001110011111101001000001001010000100010100011111010111100001001000101110011111101100101000111000010111111001100011;


module Bresenham_circle(CLOCK_50,KEY_N,SW,lockingkeyinput,vga_colour,vga_plot,vga_x,vga_y);
  input CLOCK_50;
 input [3:0] KEY_N;
 input [9:0] SW;
 input [127:0] lockingkeyinput;
 output [2:0] vga_colour;
 output vga_plot;
 output [7:0] vga_x;
 output [6:0] vga_y;
 wire _0736_;
 wire _0148_;
 wire _0619_;
 wire _0614_;
 wire _0481_;
 wire _0412_;
 wire _1035_;
 wire _0551_;
 wire _0639_;
 wire _0271_;
 wire _0623_;
 wire _0995_;
 wire _0449_;
 wire _0734_;
 wire _0345_;
 wire _0393_;
 wire _0751_;
 wire _0230_;
 wire _0097_;
 wire [7:0] T3x;
 wire _0689_;
 wire _0156_;
 wire _0849_;
 wire _0705_;
 wire _0526_;
 wire _0528_;
 wire _0073_;
 wire _0071_;
 wire _0203_;
 wire _0943_;
 wire _0452_;
 wire _0937_;
 wire _0621_;
 wire _0648_;
 wire _0740_;
 wire _0638_;
 wire _0636_;
 wire _0852_;
 wire _0173_;
 wire _0390_;
 wire _0252_;
 wire _0659_;
 wire _0598_;
 wire _0691_;
 wire _0057_;
 wire _0576_;
 wire _0758_;
 wire _0278_;
 wire _0081_;
 wire _0676_;
 wire _0229_;
 wire _0060_;
 wire _0537_;
 wire _0905_;
 wire _0202_;
 wire _0700_;
 wire _0973_;
 wire _0539_;
 wire _0624_;
 wire _0769_;
 wire _0343_;
 wire _0786_;
 wire _0075_;
 wire _0787_;
 wire _0836_;
 wire _0902_;
 wire _1020_;
 wire _0098_;
 wire _0019_;
 wire _0124_;
 wire _0126_;
 wire _0692_;
 wire _1023_;
 wire _0302_;
 wire _0738_;
 wire _0214_;
 wire _0056_;
 wire _0199_;
 wire _0702_;
 wire _0859_;
 wire _0201_;
 wire _0167_;
 wire _0867_;
 wire _0448_;
 wire _0664_;
 wire _0647_;
 wire _0851_;
 wire _0955_;
 wire _0978_;
 wire _0723_;
 wire _0674_;
 wire _0766_;
 wire _0140_;
 wire _0595_;
 wire _0105_;
 wire _0004_;
 wire _1032_;
 wire _0095_;
 wire _0086_;
 wire _1003_;
 wire _0768_;
 wire _1010_;
 wire _0834_;
 wire _0954_;
 wire _0050_;
 wire _0453_;
 wire _1026_;
 wire _0792_;
 wire _0927_;
 wire _0335_;
 wire _0036_;
 wire _0893_;
 wire _0625_;
 wire _0970_;
 wire _0891_;
 wire _0910_;
 wire _0021_;
 wire _1017_;
 wire _0361_;
 wire _0248_;
 wire _0320_;
 wire _0181_;
 wire _0699_;
 wire _0915_;
 wire _0919_;
 wire _0720_;
 wire _0532_;
 wire _0286_;
 wire _0750_;
 wire _0871_;
 wire _0498_;
 wire _0592_;
 wire _0254_;
 wire _0504_;
 wire _0832_;
 wire _0553_;
 wire _0317_;
 wire _0435_;
 wire _0548_;
 wire _0030_;
 wire _0556_;
 wire _0974_;
 wire _0425_;
 wire _0338_;
 wire _0994_;
 wire _0296_;
 wire _0487_;
 wire _0160_;
 wire _0853_;
 wire _0471_;
 wire _0022_;
 wire _0976_;
 wire _0701_;
 wire _0815_;
 wire _0318_;
 wire _0656_;
 wire _0103_;
 wire _0123_;
 wire _0336_;
 wire _0348_;
 wire _0782_;
 wire _0916_;
 wire _0074_;
 wire _0236_;
 wire _0009_;
 wire _0017_;
 wire _0039_;
 wire _0427_;
 wire _0735_;
 wire _0979_;
 wire _0277_;
 wire _0176_;
 wire _1007_;
 wire _0186_;
 wire _0323_;
 wire _0628_;
 wire _0714_;
 wire _0387_;
 wire _0831_;
 wire _0187_;
 wire _0771_;
 wire _0741_;
 wire _0847_;
 wire _0276_;
 wire _0732_;
 wire _0450_;
 wire _0053_;
 wire _0835_;
 wire _0415_;
 wire _0651_;
 wire _0055_;
 wire _0110_;
 wire _0114_;
 wire _0303_;
 wire _0262_;
 wire _0765_;
 wire _0462_;
 wire _0640_;
 wire [2:0] T3colourcircle;
 wire _1029_;
 wire _1021_;
 wire _0288_;
 wire _0465_;
 wire _0827_;
 wire _0655_;
 wire _0294_;
 wire _0228_;
 wire _0936_;
 wire _0015_;
 wire _0508_;
 wire _0145_;
 wire _0865_;
 wire _0968_;
 wire _0483_;
 wire _0096_;
 wire _0963_;
 wire _0334_;
 wire _0475_;
 wire _0028_;
 wire _0839_;
 wire _0707_;
 wire _0838_;
 wire _0856_;
 wire _0012_;
 wire _0431_;
 wire _0131_;
 wire _0143_;
 wire _1037_;
 wire _0225_;
 wire _0550_;
 wire _0562_;
 wire _0542_;
 wire _0165_;
 wire _0693_;
 wire _0660_;
 wire _0744_;
 wire _0025_;
 wire _0993_;
 wire _1014_;
 wire _0454_;
 wire _1028_;
 wire _0918_;
 wire _0269_;
 wire _0869_;
 wire _0746_;
 wire _0121_;
 wire _0668_;
 wire _0570_;
 wire _0389_;
 wire _0833_;
 wire _0613_;
 wire _0093_;
 wire _0575_;
 wire _0480_;
 wire _0468_;
 wire _0681_;
 wire _0061_;
 wire _0089_;
 wire _0312_;
 wire _0616_;
 wire _0541_;
 wire _0885_;
 wire _0281_;
 wire _0326_;
 wire _0913_;
 wire _0727_;
 wire _0533_;
 wire _0604_;
 wire _0952_;
 wire _0018_;
 wire _0185_;
 wire _0810_;
 wire _0319_;
 wire _0330_;
 wire _0922_;
 wire _0695_;
 wire _0067_;
 wire _0351_;
 wire _1016_;
 wire _0094_;
 wire _0661_;
 wire _0003_;
 wire _0384_;
 wire _0178_;
 wire _0724_;
 wire _0646_;
 wire _0710_;
 wire _0703_;
 wire _0761_;
 wire _0808_;
 wire _0799_;
 wire _0175_;
 wire _0224_;
 wire _0878_;
 wire _0418_;
 wire _0234_;
 wire _0085_;
 wire _0814_;
 wire _0423_;
 wire _0138_;
 wire _0005_;
 wire _0620_;
 wire _0256_;
 wire _0411_;
 wire _0354_;
 wire _0049_;
 wire _0408_;
 wire _0298_;
 wire T3plot;
 wire _0111_;
 wire _0293_;
 wire _0872_;
 wire _0013_;
 wire _0120_;
 wire _0109_;
 wire _0608_;
 wire _0082_;
 wire _0882_;
 wire _0581_;
 wire _0829_;
 wire _0200_;
 wire _0737_;
 wire _0823_;
 wire _0906_;
 wire _0400_;
 wire _0191_;
 wire _0797_;
 wire _0579_;
 wire _0605_;
 wire _0287_;
 wire _0934_;
 wire _0840_;
 wire _0957_;
 wire _0825_;
 wire _0899_;
 wire _0136_;
 wire _0235_;
 wire _1033_;
 wire _0374_;
 wire _0597_;
 wire _0679_;
 wire _0939_;
 wire _0554_;
 wire _0363_;
 wire _0432_;
 wire _0862_;
 wire _0622_;
 wire _0618_;
 wire _0748_;
 wire _0743_;
 wire _0889_;
 wire _0289_;
 wire _0267_;
 wire _0451_;
 wire _0297_;
 wire _0362_;
 wire _0188_;
 wire _0466_;
 wire _0985_;
 wire _0459_;
 wire _0762_;
 wire _0163_;
 wire _0924_;
 wire _0327_;
 wire _0802_;
 wire _0373_;
 wire _0244_;
 wire _0870_;
 wire _0544_;
 wire _0567_;
 wire _0458_;
 wire _0909_;
 wire _0488_;
 wire _0980_;
 wire _0369_;
 wire _0818_;
 wire _0997_;
 wire _0589_;
 wire _0784_;
 wire _0040_;
 wire _0133_;
 wire _0386_;
 wire _0329_;
 wire _1030_;
 wire _0135_;
 wire _0777_;
 wire _0255_;
 wire _0159_;
 wire _0112_;
 wire _0516_;
 wire _0938_;
 wire _0896_;
 wire _0717_;
 wire _0726_;
 wire _0972_;
 wire _0346_;
 wire _0857_;
 wire _0208_;
 wire _0195_;
 wire _0383_;
 wire _0099_;
 wire _0530_;
 wire _0520_;
 wire _0880_;
 wire _0051_;
 wire _0804_;
 wire _0926_;
 wire _0014_;
 wire _0440_;
 wire _0557_;
 wire _1024_;
 wire _0394_;
 wire _0945_;
 wire _0967_;
 wire _0713_;
 wire _0593_;
 wire _0990_;
 wire _0032_;
 wire _0037_;
 wire _0983_;
 wire _0006_;
 wire _0630_;
 wire _0644_;
 wire _0301_;
 wire _0884_;
 wire _0992_;
 wire _0194_;
 wire _0842_;
 wire _0642_;
 wire _0645_;
 wire _0672_;
 wire _0966_;
 wire _0058_;
 wire _0359_;
 wire _0401_;
 wire _0333_;
 wire _0908_;
 wire _0812_;
 wire _0391_;
 wire _0753_;
 wire _0137_;
 wire _0629_;
 wire _0845_;
 wire _1015_;
 wire _0986_;
 wire _0091_;
 wire _0356_;
 wire _0168_;
 wire _0684_;
 wire _0026_;
 wire _0344_;
 wire _0685_;
 wire _0065_;
 wire _0903_;
 wire _0023_;
 wire [2:0] T2colour;
 wire _0162_;
 wire _0239_;
 wire _0113_;
 wire _0883_;
 wire _0282_;
 wire _0848_;
 wire _0935_;
 wire _0585_;
 wire _0694_;
 wire _0339_;
 wire _0396_;
 wire _0868_;
 wire _1001_;
 wire _0456_;
 wire _0873_;
 wire _0180_;
 wire _0237_;
 wire _0001_;
 wire _0545_;
 wire _0147_;
 wire _0219_;
 wire _0590_;
 wire _0261_;
 wire _0923_;
 wire _1012_;
 wire _0901_;
 wire _0414_;
 wire _1027_;
 wire _0441_;
 wire _0424_;
 wire _0409_;
 wire _0158_;
 wire _0007_;
 wire _0772_;
 wire _0300_;
 wire _0874_;
 wire _0779_;
 wire _0259_;
 wire _0042_;
 wire _0117_;
 wire _0569_;
 wire _1009_;
 wire _0217_;
 wire _0951_;
 wire _0206_;
 wire _0855_;
 wire _1000_;
 wire _0665_;
 wire _0828_;
 wire _0041_;
 wire _0875_;
 wire _0864_;
 wire _0601_;
 wire _0977_;
 wire _0637_;
 wire _0139_;
 wire [6:0] T3yp;
 wire _0299_;
 wire _0008_;
 wire _0045_;
 wire _0603_;
 wire _0382_;
 wire _0775_;
 wire _0912_;
 wire _0580_;
 wire _0315_;
 wire _0207_;
 wire _0560_;
 wire _0170_;
 wire _0034_;
 wire _0552_;
 wire _0398_;
 wire _0730_;
 wire _0144_;
 wire _0523_;
 wire _0104_;
 wire _0770_;
 wire _0555_;
 wire _0245_;
 wire _0265_;
 wire _0474_;
 wire _0166_;
 wire _0249_;
 wire _0410_;
 wire _0273_;
 wire _0756_;
 wire _0337_;
 wire _0325_;
 wire _0843_;
 wire _0958_;
 wire _0830_;
 wire _0760_;
 wire _0960_;
 wire _0381_;
 wire _0931_;
 wire _0485_;
 wire _0650_;
 wire _0774_;
 wire _0024_;
 wire _0634_;
 wire _0793_;
 wire _0538_;
 wire _0503_;
 wire _0584_;
 wire _0610_;
 wire _0984_;
 wire _0791_;
 wire _0029_;
 wire _0090_;
 wire _0063_;
 wire _0500_;
 wire _0698_;
 wire _0472_;
 wire _1019_;
 wire _0101_;
 wire _0632_;
 wire _0031_;
 wire _0591_;
 wire _0989_;
 wire _0011_;
 wire T2Done;
 wire _0725_;
 wire _0118_;
 wire [7:0] T3xp;
 wire _1036_;
 wire _1025_;
 wire _0275_;
 wire _0971_;
 wire _0182_;
 wire _0146_;
 wire _0800_;
 wire _0129_;
 wire _0446_;
 wire _0921_;
 wire _0429_;
 wire _0861_;
 wire _0745_;
 wire _0434_;
 wire _0284_;
 wire _0780_;
 wire _1008_;
 wire _0502_;
 wire _0559_;
 wire _0246_;
 wire _0455_;
 wire _0377_;
 wire _0379_;
 wire _0494_;
 wire _0731_;
 wire _0649_;
 wire _0107_;
 wire _0308_;
 wire _0981_;
 wire _0179_;
 wire _0305_;
 wire _0953_;
 wire _0657_;
 wire _0413_;
 wire _0663_;
 wire _0263_;
 wire _0611_;
 wire _0033_;
 wire _0606_;
 wire _0406_;
 wire _0577_;
 wire _1004_;
 wire _0524_;
 wire _0654_;
 wire _0285_;
 wire _0493_;
 wire _0238_;
 wire _0052_;
 wire _0599_;
 wire _0368_;
 wire _0566_;
 wire _0304_;
 wire _0059_;
 wire _0515_;
 wire _0749_;
 wire _0347_;
 wire _0438_;
 wire _0397_;
 wire _0077_;
 wire _0227_;
 wire _0422_;
 wire _0242_;
 wire _1011_;
 wire _0027_;
 wire _0641_;
 wire _0820_;
 wire _0380_;
 wire _0948_;
 wire _0084_;
 wire _0546_;
 wire _0243_;
 wire _0813_;
 wire _0805_;
 wire _0711_;
 wire _0962_;
 wire _0739_;
 wire _0505_;
 wire _0106_;
 wire _0959_;
 wire _1022_;
 wire _0688_;
 wire _0988_;
 wire _0100_;
 wire _0080_;
 wire _0788_;
 wire _0911_;
 wire _0416_;
 wire _0907_;
 wire _0247_;
 wire _0667_;
 wire _1034_;
 wire _0125_;
 wire _0222_;
 wire _0274_;
 wire _0587_;
 wire _0314_;
 wire _0757_;
 wire _0122_;
 wire _0858_;
 wire _0460_;
 wire _0241_;
 wire _0671_;
 wire _0342_;
 wire _0961_;
 wire _0690_;
 wire T2plot;
 wire _0189_;
 wire _0817_;
 wire _0436_;
 wire _0897_;
 wire _0283_;
 wire _0933_;
 wire _0421_;
 wire _0594_;
 wire _0212_;
 wire _0819_;
 wire _0811_;
 wire _0469_;
 wire _0445_;
 wire _0047_;
 wire _0439_;
 wire _0164_;
 wire _0280_;
 wire _0941_;
 wire _1006_;
 wire _0708_;
 wire _0038_;
 wire _1018_;
 wire _0627_;
 wire _0108_;
 wire _0824_;
 wire _0999_;
 wire _0192_;
 wire _0420_;
 wire _0841_;
 wire _0549_;
 wire _0742_;
 wire _0444_;
 wire _0064_;
 wire _0678_;
 wire _0221_;
 wire _0816_;
 wire _0115_;
 wire _0430_;
 wire _0783_;
 wire _0132_;
 wire _0716_;
 wire _0352_;
 wire _0291_;
 wire _0615_;
 wire _0733_;
 wire _0251_;
 wire _0322_;
 wire _0572_;
 wire _0881_;
 wire _0403_;
 wire _0950_;
 wire _0232_;
 wire _0582_;
 wire _1031_;
 wire _0174_;
 wire _0177_;
 wire _0917_;
 wire _0321_;
 wire _0443_;
 wire _0586_;
 wire _0155_;
 wire _0171_;
 wire _0290_;
 wire _0470_;
 wire _0510_;
 wire _0790_;
 wire _0169_;
 wire _0371_;
 wire _0876_;
 wire _0602_;
 wire _0204_;
 wire _0925_;
 wire _0486_;
 wire _0358_;
 wire _0998_;
 wire _0193_;
 wire _0670_;
 wire _0755_;
 wire [3:0] T3state;
 wire _0044_;
 wire _0332_;
 wire _0509_;
 wire _0519_;
 wire _0484_;
 wire _0696_;
 wire _0066_;
 wire _0153_;
 wire _0571_;
 wire _0512_;
 wire _0464_;
 wire _0404_;
 wire _0257_;
 wire _0877_;
 wire _0956_;
 wire _0209_;
 wire _0054_;
 wire _0965_;
 wire _0324_;
 wire _0392_;
 wire _0079_;
 wire _0215_;
 wire _0405_;
 wire _0152_;
 wire _0331_;
 wire _0540_;
 wire _0767_;
 wire _0130_;
 wire _0525_;
 wire _0890_;
 wire _0355_;
 wire _0798_;
 wire _0437_;
 wire _0478_;
 wire _0310_;
 wire _0399_;
 wire _0428_;
 wire _0596_;
 wire _0272_;
 wire _0653_;
 wire _0360_;
 wire _0850_;
 wire _0072_;
 wire _0020_;
 wire _0666_;
 wire _0947_;
 wire _0076_;
 wire _0534_;
 wire _0506_;
 wire _0673_;
 wire _0035_;
 wire _0803_;
 wire _0609_;
 wire _0489_;
 wire _0491_;
 wire _0987_;
 wire _0309_;
 wire _0365_;
 wire _0311_;
 wire _0894_;
 wire _0388_;
 wire _0776_;
 wire _0914_;
 wire _0643_;
 wire _0563_;
 wire _0497_;
 wire _0417_;
 wire _0573_;
 wire _0975_;
 wire _1013_;
 wire _0376_;
 wire _0709_;
 wire _0395_;
 wire _0796_;
 wire _0226_;
 wire _0795_;
 wire _0617_;
 wire _0016_;
 wire _0531_;
 wire _0759_;
 wire _0892_;
 wire _0461_;
 wire _0102_;
 wire _0529_;
 wire _0535_;
 wire _0205_;
 wire _0270_;
 wire _0801_;
 wire _0295_;
 wire _0198_;
 wire _0141_;
 wire _0210_;
 wire _0433_;
 wire _0754_;
 wire _0157_;
 wire _0340_;
 wire _0558_;
 wire _0860_;
 wire _0518_;
 wire _0378_;
 wire _0062_;
 wire _0316_;
 wire _0088_;
 wire _0353_;
 wire _0341_;
 wire _0069_;
 wire _0982_;
 wire _0887_;
 wire _0197_;
 wire _0048_;
 wire _0211_;
 wire _0949_;
 wire _0279_;
 wire _0231_;
 wire _0092_;
 wire _0149_;
 wire _0266_;
 wire _0942_;
 wire _0564_;
 wire _0264_;
 wire _0675_;
 wire _0511_;
 wire _0600_;
 wire _0729_;
 wire _0514_;
 wire _0578_;
 wire _0932_;
 wire _0495_;
 wire _0078_;
 wire _0807_;
 wire _0522_;
 wire _0929_;
 wire _0292_;
 wire _0366_;
 wire _0728_;
 wire _0463_;
 wire _0879_;
 wire _0083_;
 wire _0499_;
 wire _0151_;
 wire _0677_;
 wire _0161_;
 wire _0612_;
 wire _0778_;
 wire _0043_;
 wire _1002_;
 wire _0184_;
 wire _0658_;
 wire _0996_;
 wire _0119_;
 wire _0821_;
 wire _0631_;
 wire _0719_;
 wire _0822_;
 wire _0220_;
 wire _0863_;
 wire _0240_;
 wire _0442_;
 wire _0476_;
 wire _0218_;
 wire _0785_;
 wire _0898_;
 wire _0154_;
 wire _0070_;
 wire _0258_;
 wire _0457_;
 wire _0196_;
 wire _0763_;
 wire [7:0] T2x;
 wire _0002_;
 wire _0928_;
 wire _0633_;
 wire _0930_;
 wire _0781_;
 wire _0991_;
 wire _0568_;
 wire _0652_;
 wire _0473_;
 wire _0715_;
 wire _0826_;
 wire _0547_;
 wire _0794_;
 wire [8:0] T3d;
 wire _0507_;
 wire _0357_;
 wire _0944_;
 wire _0704_;
 wire _0752_;
 wire _0895_;
 wire _0127_;
 wire _0964_;
 wire _0313_;
 wire _0721_;
 wire _0583_;
 wire _0722_;
 wire _0946_;
 wire _0367_;
 wire _0536_;
 wire _0588_;
 wire _0306_;
 wire _0350_;
 wire _0407_;
 wire _0940_;
 wire _0626_;
 wire _0134_;
 wire _0087_;
 wire _0496_;
 wire _0477_;
 wire _0517_;
 wire _0682_;
 wire _0662_;
 wire _0128_;
 wire _0846_;
 wire _0068_;
 wire _0886_;
 wire _0706_;
 wire _0969_;
 wire _0686_;
 wire _0635_;
 wire _0233_;
 wire _0213_;
 wire _0490_;
 wire _0190_;
 wire _0402_;
 wire _0513_;
 wire _0561_;
 wire _0010_;
 wire _0574_;
 wire _0000_;
 wire _0565_;
 wire _0764_;
 wire _0866_;
 wire _0501_;
 wire _0253_;
 wire _0223_;
 wire _0904_;
 wire _0328_;
 wire _0669_;
 wire _0046_;
 wire _0888_;
 wire _0419_;
 wire _0150_;
 wire _0920_;
 wire _0900_;
 wire _0307_;
 wire _0385_;
 wire _0773_;
 wire _0747_;
 wire _0447_;
 wire [6:0] T3y;
 wire _0250_;
 wire _0844_;
 wire _0375_;
 wire _0809_;
 wire _0260_;
 wire _0172_;
 wire _0492_;
 wire _0543_;
 wire _0521_;
 wire _0370_;
 wire _0837_;
 wire _0482_;
 wire _0216_;
 wire _0607_;
 wire _0372_;
 wire _0467_;
 wire _1005_;
 wire _0426_;
 wire _0712_;
 wire _0854_;
 wire _0349_;
 wire _0697_;
 wire _0789_;
 wire _0364_;
 wire _0268_;
 wire _0183_;
 wire _0527_;
 wire _0680_;
 wire _0806_;
 wire _0479_;
 wire [6:0] T2y;
 wire _0683_;
 wire _0718_;
 wire _0687_;
 wire _0142_;
 wire _0116_;
 wire keywire1051;
 wire keywire1052;
 wire keywire1053;
 wire keywire1054;
 wire keywire1055;
 wire keywire1056;
 wire keywire1057;
 wire keywire1058;
 wire keywire1059;
 wire keywire1060;
 wire keywire1061;
 wire keywire1062;
 wire keywire1063;
 wire keywire1064;
 wire keywire1065;
 wire keywire1066;
 wire keywire1067;
 wire keywire1068;
 wire keywire1069;
 wire keywire1070;
 wire keywire1071;
 wire keywire1072;
 wire keywire1073;
 wire keywire1074;
 wire keywire1075;
 wire keywire1076;
 wire keywire1077;
 wire keywire1078;
 wire keywire1079;
 wire keywire1080;
 wire keywire1081;
 wire keywire1082;
 wire keywire1083;
 wire keywire1084;
 wire keywire1085;
 wire keywire1086;
 wire keywire1087;
 wire keywire1088;
 wire keywire1089;
 wire keywire1090;
 wire keywire1091;
 wire keywire1092;
 wire keywire1093;
 wire keywire1094;
 wire keywire1095;
 wire keywire1096;
 wire keywire1097;
 wire keywire1098;
 wire keywire1099;
 wire keywire1100;
 wire keywire1101;
 wire keywire1102;
 wire keywire1103;
 wire keywire1104;
 wire keywire1105;
 wire keywire1106;
 wire keywire1107;
 wire keywire1108;
 wire keywire1109;
 wire keywire1110;
 wire keywire1111;
 wire keywire1112;
 wire keywire1113;
 wire keywire1114;
 wire keywire1115;
 wire keywire1116;
 wire keywire1117;
 wire keywire1118;
 wire keywire1119;
 wire keywire1120;
 wire keywire1121;
 wire keywire1122;
 wire keywire1123;
 wire keywire1124;
 wire keywire1125;
 wire keywire1126;
 wire keywire1127;
 wire keywire1128;
 wire keywire1129;
 wire keywire1130;
 wire keywire1131;
 wire keywire1132;
 wire keywire1133;
 wire keywire1134;
 wire keywire1135;
 wire keywire1136;
 wire keywire1137;
 wire keywire1138;
 wire keywire1139;
 wire keywire1140;
 wire keywire1141;
 wire keywire1142;
 wire keywire1143;
 wire keywire1144;
 wire keywire1145;
 wire keywire1146;
 wire keywire1147;
 wire keywire1148;
 wire keywire1149;
 wire keywire1150;
 wire keywire1151;
 wire keywire1152;
 wire keywire1153;
 wire keywire1154;
 wire keywire1155;
 wire keywire1156;
 wire keywire1157;
 wire keywire1158;
 wire keywire1159;
 wire keywire1160;
 wire keywire1161;
 wire keywire1162;
 wire keywire1163;
 wire keywire1164;
 wire keywire1165;
 wire keywire1166;
 wire keywire1167;
 wire keywire1168;
 wire keywire1169;
 wire keywire1170;
 wire keywire1171;
 wire keywire1172;
 wire keywire1173;
 wire keywire1174;
 wire keywire1175;
 wire keywire1176;
 wire keywire1177;
 wire keywire1178;
 NOT_g NOT_1038_(.A(T2Done), .Y(_0011_));
 NOT_g NOT_1096_(.A(T2y[0]), .Y(_0113_));
 NOT_g NOT_1097_(.A(_0039_), .Y(T2plot));
 NOT_g NOT_1098_(.A(T2x[7]), .Y(keywire1177));
 NOT_g NOT_1099_(.A(T2x[6]), .Y(keywire1173));
 NOT_g NOT_1100_(.A(KEY_N[3]), .Y(keywire1118));
 NOT_g NOT_1156_(.A(_0088_), .Y(_0089_));
 NOT_g NOT_1191_(.A(KEY_N[3]), .Y(keywire1119));
 NOT_g NOT_1192_(.A(KEY_N[3]), .Y(keywire1120));
 NOT_g NOT_1193_(.A(KEY_N[3]), .Y(keywire1121));
 NOT_g NOT_1194_(.A(KEY_N[3]), .Y(keywire1122));
 NOT_g NOT_1195_(.A(KEY_N[3]), .Y(keywire1123));
 NOT_g NOT_1196_(.A(KEY_N[3]), .Y(keywire1124));
 NOT_g NOT_1197_(.A(KEY_N[3]), .Y(keywire1125));
 NOT_g NOT_1198_(.A(KEY_N[3]), .Y(keywire1126));
 NOT_g NOT_1199_(.A(KEY_N[3]), .Y(keywire1127));
 NOT_g NOT_1200_(.A(KEY_N[3]), .Y(keywire1128));
 NOT_g NOT_1201_(.A(KEY_N[3]), .Y(keywire1129));
 NOT_g NOT_1202_(.A(KEY_N[3]), .Y(keywire1130));
 NOT_g NOT_1203_(.A(KEY_N[3]), .Y(keywire1131));
 NOT_g NOT_1204_(.A(KEY_N[3]), .Y(keywire1132));
 NOT_g NOT_1205_(.A(KEY_N[3]), .Y(keywire1133));
 NOT_g NOT_1226_(.A(T3state[3]), .Y(_0210_));
 NOT_g NOT_1227_(.A(T3state[2]), .Y(_0211_));
 NOT_g NOT_1228_(.A(T3state[0]), .Y(_0212_));
 NOT_g NOT_1229_(.A(KEY_N[3]), .Y(keywire1134));
 NOT_g NOT_1230_(.A(T3y[0]), .Y(_0213_));
 NOT_g NOT_1231_(.A(T3y[1]), .Y(_0214_));
 NOT_g NOT_1232_(.A(T3y[2]), .Y(_0215_));
 NOT_g NOT_1233_(.A(T3y[3]), .Y(_0216_));
 NOT_g NOT_1234_(.A(T3y[4]), .Y(_0217_));
 NOT_g NOT_1235_(.A(T3y[5]), .Y(_0218_));
 NOT_g NOT_1236_(.A(T3y[6]), .Y(_0219_));
 NOT_g NOT_1237_(.A(T3d[1]), .Y(_0220_));
 NOT_g NOT_1238_(.A(T3x[0]), .Y(_0221_));
 NOT_g NOT_1239_(.A(T3x[1]), .Y(_0222_));
 NOT_g NOT_1240_(.A(T3x[2]), .Y(_0223_));
 NOT_g NOT_1241_(.A(T3x[3]), .Y(_0224_));
 NOT_g NOT_1242_(.A(T3x[4]), .Y(_0225_));
 NOT_g NOT_1243_(.A(T3x[5]), .Y(_0226_));
 NOT_g NOT_1244_(.A(T3x[6]), .Y(_0227_));
 NOT_g NOT_1245_(.A(SW[3]), .Y(keywire1142));
 NOT_g NOT_1246_(.A(SW[4]), .Y(keywire1143));
 NOT_g NOT_1247_(.A(1'h1), .Y(_0230_));
 NOT_g NOT_1248_(.A(1'h1), .Y(_0231_));
 NOT_g NOT_1249_(.A(1'h0), .Y(_0232_));
 NOT_g NOT_1250_(.A(1'h1), .Y(_0233_));
 NOT_g NOT_1251_(.A(1'h1), .Y(_0234_));
 NOT_g NOT_1252_(.A(1'h1), .Y(_0235_));
 NOT_g NOT_1262_(.A(_0244_), .Y(_0245_));
 NOT_g NOT_1266_(.A(_0248_), .Y(_0249_));
 NOT_g NOT_1270_(.A(_0252_), .Y(_0253_));
 NOT_g NOT_1322_(.A(_0301_), .Y(T3plot));
 NOT_g NOT_1341_(.A(_0318_), .Y(_0319_));
 NOT_g NOT_1359_(.A(_0335_), .Y(_0336_));
 NOT_g NOT_1407_(.A(_0374_), .Y(_0375_));
 NOT_g NOT_1645_(.A(_0604_), .Y(_0175_));
 NOT_g NOT_1721_(.A(_0676_), .Y(_0677_));
 NOT_g NOT_1785_(.A(_0738_), .Y(_0739_));
 NOT_g NOT_1969_(.A(_0908_), .Y(_0909_));
 NOT_g NOT_1972_(.A(_0911_), .Y(_0912_));
 NOT_g NOT_1982_(.A(_0921_), .Y(_0922_));
 NOT_g NOT_1985_(.A(_0924_), .Y(_0925_));
 NOT_g NOT_2113_(.A(KEY_N[3]), .Y(keywire1135));
 NOT_g NOT_2114_(.A(KEY_N[3]), .Y(keywire1136));
 NOT_g NOT_2115_(.A(KEY_N[3]), .Y(keywire1137));
 NAND_g NAND_1039_(.A(T2Done), .B(T3colourcircle[0]), .Y(_0012_));
 NAND_g NAND_1040_(.A(_0011_), .B(T2colour[0]), .Y(_0013_));
 NAND_g NAND_1041_(.A(_0013_), .B(_0012_), .Y(vga_colour[0]));
 NAND_g NAND_1042_(.A(T3colourcircle[1]), .B(T2Done), .Y(_0014_));
 NAND_g NAND_1043_(.A(T2colour[1]), .B(_0011_), .Y(_0015_));
 NAND_g NAND_1044_(.A(_0015_), .B(_0014_), .Y(vga_colour[1]));
 NAND_g NAND_1045_(.A(T3colourcircle[2]), .B(T2Done), .Y(_0016_));
 NAND_g NAND_1046_(.A(T2colour[2]), .B(_0011_), .Y(_0017_));
 NAND_g NAND_1047_(.A(_0017_), .B(_0016_), .Y(vga_colour[2]));
 NAND_g NAND_1048_(.A(T3plot), .B(T2Done), .Y(_0018_));
 NAND_g NAND_1049_(.A(T2plot), .B(_0011_), .Y(_0019_));
 NAND_g NAND_1050_(.A(_0019_), .B(_0018_), .Y(vga_plot));
 NAND_g NAND_1051_(.A(T3yp[0]), .B(T2Done), .Y(_0020_));
 NAND_g NAND_1052_(.A(T2y[0]), .B(_0011_), .Y(_0021_));
 NAND_g NAND_1053_(.A(_0021_), .B(_0020_), .Y(vga_y[0]));
 NAND_g NAND_1054_(.A(T3yp[1]), .B(T2Done), .Y(_0022_));
 NAND_g NAND_1055_(.A(T2y[1]), .B(_0011_), .Y(_0023_));
 NAND_g NAND_1056_(.A(_0023_), .B(_0022_), .Y(vga_y[1]));
 NAND_g NAND_1057_(.A(T3yp[2]), .B(T2Done), .Y(_0024_));
 NAND_g NAND_1058_(.A(T2y[2]), .B(_0011_), .Y(_0025_));
 NAND_g NAND_1059_(.A(_0025_), .B(_0024_), .Y(vga_y[2]));
 NAND_g NAND_1060_(.A(T3yp[3]), .B(T2Done), .Y(_0026_));
 NAND_g NAND_1061_(.A(T2y[3]), .B(_0011_), .Y(_0027_));
 NAND_g NAND_1062_(.A(_0027_), .B(_0026_), .Y(vga_y[3]));
 NAND_g NAND_1063_(.A(T3yp[4]), .B(T2Done), .Y(_0028_));
 NAND_g NAND_1064_(.A(T2y[4]), .B(_0011_), .Y(_0029_));
 NAND_g NAND_1065_(.A(_0029_), .B(_0028_), .Y(vga_y[4]));
 NAND_g NAND_1066_(.A(T3yp[5]), .B(T2Done), .Y(_0030_));
 NAND_g NAND_1067_(.A(T2y[5]), .B(_0011_), .Y(_0031_));
 NAND_g NAND_1068_(.A(_0031_), .B(_0030_), .Y(vga_y[5]));
 NAND_g NAND_1069_(.A(T3yp[6]), .B(T2Done), .Y(_0032_));
 NAND_g NAND_1070_(.A(T2y[6]), .B(_0011_), .Y(_0033_));
 NAND_g NAND_1071_(.A(_0033_), .B(_0032_), .Y(vga_y[6]));
 NAND_g NAND_1072_(.A(T3xp[0]), .B(T2Done), .Y(_0034_));
 NAND_g NAND_1073_(.A(T2x[0]), .B(_0011_), .Y(keywire1155));
 NAND_g NAND_1074_(.A(_0035_), .B(_0034_), .Y(vga_x[0]));
 NAND_g NAND_1075_(.A(T3xp[1]), .B(T2Done), .Y(_0036_));
 NAND_g NAND_1076_(.A(T2x[1]), .B(_0011_), .Y(keywire1159));
 NAND_g NAND_1077_(.A(_0037_), .B(_0036_), .Y(vga_x[1]));
 NAND_g NAND_1078_(.A(T3xp[2]), .B(T2Done), .Y(_0038_));
 NAND_g NAND_1079_(.A(T2x[2]), .B(_0011_), .Y(keywire1160));
 NAND_g NAND_1080_(.A(_0000_), .B(_0038_), .Y(vga_x[2]));
 NAND_g NAND_1081_(.A(T3xp[3]), .B(T2Done), .Y(_0001_));
 NAND_g NAND_1082_(.A(T2x[3]), .B(_0011_), .Y(keywire1163));
 NAND_g NAND_1083_(.A(_0002_), .B(_0001_), .Y(vga_x[3]));
 NAND_g NAND_1084_(.A(T3xp[4]), .B(T2Done), .Y(_0003_));
 NAND_g NAND_1085_(.A(T2x[4]), .B(_0011_), .Y(keywire1166));
 NAND_g NAND_1086_(.A(_0004_), .B(_0003_), .Y(vga_x[4]));
 NAND_g NAND_1087_(.A(T3xp[5]), .B(T2Done), .Y(_0005_));
 NAND_g NAND_1088_(.A(T2x[5]), .B(_0011_), .Y(keywire1169));
 NAND_g NAND_1089_(.A(_0006_), .B(_0005_), .Y(keywire1051));
 NAND_g NAND_1090_(.A(T3xp[6]), .B(T2Done), .Y(_0007_));
 NAND_g NAND_1091_(.A(T2x[6]), .B(_0011_), .Y(keywire1174));
 NAND_g NAND_1092_(.A(_0008_), .B(_0007_), .Y(vga_x[6]));
 NAND_g NAND_1093_(.A(T3xp[7]), .B(T2Done), .Y(_0009_));
 NAND_g NAND_1094_(.A(T2x[7]), .B(_0011_), .Y(keywire1178));
 NAND_g NAND_1095_(.A(_0010_), .B(_0009_), .Y(vga_x[7]));
 NAND_g NAND_1108_(.A(_0121_), .B(_0119_), .Y(_0123_));
 NAND_g NAND_1112_(.A(_0126_), .B(T2y[4]), .Y(_0127_));
 NAND_g NAND_1115_(.A(_0129_), .B(_0122_), .Y(_0130_));
 NAND_g NAND_1116_(.A(_0130_), .B(T2plot), .Y(_0071_));
 NAND_g NAND_1124_(.A(_0137_), .B(_0115_), .Y(_0138_));
 NAND_g NAND_1126_(.A(_0138_), .B(T2x[7]), .Y(_0140_));
 NAND_g NAND_1127_(.A(_0139_), .B(_0130_), .Y(_0141_));
 NAND_g NAND_1132_(.A(_0141_), .B(T2y[5]), .Y(_0145_));
 NAND_g NAND_1134_(.A(_0146_), .B(_0133_), .Y(_0147_));
 NAND_g NAND_1135_(.A(_0147_), .B(_0145_), .Y(_0069_));
 NAND_g NAND_1136_(.A(_0141_), .B(T2y[4]), .Y(_0148_));
 NAND_g NAND_1138_(.A(_0075_), .B(_0133_), .Y(_0076_));
 NAND_g NAND_1139_(.A(_0076_), .B(_0148_), .Y(_0068_));
 NAND_g NAND_1140_(.A(_0140_), .B(T2y[3]), .Y(_0077_));
 NAND_g NAND_1142_(.A(_0078_), .B(_0133_), .Y(_0079_));
 NAND_g NAND_1143_(.A(_0079_), .B(_0077_), .Y(_0067_));
 NAND_g NAND_1144_(.A(_0141_), .B(T2y[2]), .Y(_0080_));
 NAND_g NAND_1146_(.A(_0081_), .B(_0133_), .Y(_0082_));
 NAND_g NAND_1147_(.A(_0082_), .B(_0080_), .Y(_0066_));
 NAND_g NAND_1148_(.A(_0141_), .B(T2y[1]), .Y(_0083_));
 NAND_g NAND_1150_(.A(_0084_), .B(_0133_), .Y(_0085_));
 NAND_g NAND_1151_(.A(_0085_), .B(_0083_), .Y(_0065_));
 NAND_g NAND_1152_(.A(_0133_), .B(_0113_), .Y(_0086_));
 NAND_g NAND_1153_(.A(_0141_), .B(T2y[0]), .Y(_0087_));
 NAND_g NAND_1154_(.A(_0087_), .B(_0086_), .Y(_0064_));
 NAND_g NAND_1157_(.A(_0088_), .B(T2x[6]), .Y(keywire1175));
 NAND_g NAND_1158_(.A(_0090_), .B(_0114_), .Y(_0091_));
 NAND_g NAND_1165_(.A(_0094_), .B(_0140_), .Y(_0095_));
 NAND_g NAND_1166_(.A(_0095_), .B(_0130_), .Y(_0060_));
 NAND_g NAND_1168_(.A(_0096_), .B(_0140_), .Y(_0097_));
 NAND_g NAND_1169_(.A(_0097_), .B(_0130_), .Y(_0059_));
 NAND_g NAND_1171_(.A(_0098_), .B(_0140_), .Y(_0099_));
 NAND_g NAND_1172_(.A(_0099_), .B(_0130_), .Y(_0058_));
 NAND_g NAND_1174_(.A(_0100_), .B(_0140_), .Y(_0101_));
 NAND_g NAND_1175_(.A(_0101_), .B(_0130_), .Y(_0057_));
 NAND_g NAND_1176_(.A(_0130_), .B(T2x[0]), .Y(keywire1156));
 NAND_g NAND_1179_(.A(T2y[0]), .B(SW[9]), .Y(keywire1152));
 NAND_g NAND_1183_(.A(T2y[1]), .B(SW[9]), .Y(keywire1153));
 NAND_g NAND_1187_(.A(SW[9]), .B(T2y[2]), .Y(keywire1154));
 NAND_g NAND_1255_(.A(_0236_), .B(_0211_), .Y(_0238_));
 NAND_g NAND_1257_(.A(_0238_), .B(T3state[3]), .Y(_0240_));
 NAND_g NAND_1259_(.A(_0240_), .B(T2Done), .Y(_0242_));
 NAND_g NAND_1261_(.A(_0243_), .B(_0215_), .Y(_0244_));
 NAND_g NAND_1265_(.A(_0247_), .B(_0218_), .Y(_0248_));
 NAND_g NAND_1271_(.A(_0252_), .B(T3state[1]), .Y(_0254_));
 NAND_g NAND_1276_(.A(_0251_), .B(_0236_), .Y(_0258_));
 NAND_g NAND_1279_(.A(_0260_), .B(T3state[1]), .Y(_0261_));
 NAND_g NAND_1280_(.A(_0261_), .B(_0258_), .Y(_0262_));
 NAND_g NAND_1285_(.A(_0242_), .B(_0211_), .Y(_0267_));
 NAND_g NAND_1286_(.A(_0266_), .B(_0241_), .Y(_0268_));
 NAND_g NAND_1288_(.A(_0242_), .B(T3state[1]), .Y(_0269_));
 NAND_g NAND_1290_(.A(_0270_), .B(_0210_), .Y(_0271_));
 NAND_g NAND_1291_(.A(_0271_), .B(_0269_), .Y(_0154_));
 NAND_g NAND_1292_(.A(_0227_), .B(T3y[6]), .Y(_0272_));
 NAND_g NAND_1293_(.A(T3x[5]), .B(_0218_), .Y(_0273_));
 NAND_g NAND_1294_(.A(_0224_), .B(T3y[3]), .Y(_0274_));
 NAND_g NAND_1295_(.A(T3x[2]), .B(_0215_), .Y(_0275_));
 NAND_g NAND_1296_(.A(T3x[1]), .B(_0214_), .Y(_0276_));
 NAND_g NAND_1297_(.A(T3x[0]), .B(_0213_), .Y(_0277_));
 NAND_g NAND_1298_(.A(_0277_), .B(_0276_), .Y(_0278_));
 NAND_g NAND_1299_(.A(_0222_), .B(T3y[1]), .Y(_0279_));
 NAND_g NAND_1300_(.A(_0223_), .B(T3y[2]), .Y(_0280_));
 NAND_g NAND_1302_(.A(_0281_), .B(_0278_), .Y(_0282_));
 NAND_g NAND_1303_(.A(_0282_), .B(_0275_), .Y(_0283_));
 NAND_g NAND_1304_(.A(_0283_), .B(_0274_), .Y(_0284_));
 NAND_g NAND_1305_(.A(T3x[4]), .B(_0217_), .Y(_0285_));
 NAND_g NAND_1306_(.A(T3x[3]), .B(_0216_), .Y(_0286_));
 NAND_g NAND_1308_(.A(_0287_), .B(_0284_), .Y(_0288_));
 NAND_g NAND_1309_(.A(_0226_), .B(T3y[5]), .Y(_0289_));
 NAND_g NAND_1310_(.A(_0225_), .B(T3y[4]), .Y(_0290_));
 NAND_g NAND_1312_(.A(_0291_), .B(_0288_), .Y(_0292_));
 NAND_g NAND_1313_(.A(_0292_), .B(_0273_), .Y(_0293_));
 NAND_g NAND_1314_(.A(_0293_), .B(_0272_), .Y(_0294_));
 NAND_g NAND_1316_(.A(_0237_), .B(T3state[3]), .Y(_0296_));
 NAND_g NAND_1318_(.A(T3x[6]), .B(_0219_), .Y(_0298_));
 NAND_g NAND_1320_(.A(_0299_), .B(_0294_), .Y(_0300_));
 NAND_g NAND_1324_(.A(_0263_), .B(_0251_), .Y(_0303_));
 NAND_g NAND_1325_(.A(_0263_), .B(_0259_), .Y(_0304_));
 NAND_g NAND_1326_(.A(_0304_), .B(_0258_), .Y(_0305_));
 NAND_g NAND_1329_(.A(_0307_), .B(_0300_), .Y(_0308_));
 NAND_g NAND_1330_(.A(_0308_), .B(_0241_), .Y(_0309_));
 NAND_g NAND_1331_(.A(_0242_), .B(T3state[0]), .Y(_0310_));
 NAND_g NAND_1332_(.A(_0310_), .B(_0309_), .Y(_0153_));
 NAND_g NAND_1339_(.A(_0316_), .B(_0313_), .Y(_0317_));
 NAND_g NAND_1340_(.A(_0317_), .B(T3d[8]), .Y(_0318_));
 NAND_g NAND_1344_(.A(_0321_), .B(T3y[0]), .Y(_0322_));
 NAND_g NAND_1347_(.A(_0324_), .B(_0323_), .Y(_0325_));
 NAND_g NAND_1353_(.A(_0330_), .B(_0322_), .Y(_0157_));
 NAND_g NAND_1354_(.A(_0321_), .B(T3y[1]), .Y(_0331_));
 NAND_g NAND_1356_(.A(_0332_), .B(_0328_), .Y(_0333_));
 NAND_g NAND_1357_(.A(_0325_), .B(_0229_), .Y(_0334_));
 NAND_g NAND_1358_(.A(_0334_), .B(_0301_), .Y(_0335_));
 NAND_g NAND_1361_(.A(_0337_), .B(_0331_), .Y(_0158_));
 NAND_g NAND_1362_(.A(_0320_), .B(_0243_), .Y(_0338_));
 NAND_g NAND_1364_(.A(_0339_), .B(_0338_), .Y(_0340_));
 NAND_g NAND_1367_(.A(_0341_), .B(_0325_), .Y(_0343_));
 NAND_g NAND_1368_(.A(_0328_), .B(_0245_), .Y(_0344_));
 NAND_g NAND_1370_(.A(_0345_), .B(_0340_), .Y(_0159_));
 NAND_g NAND_1371_(.A(_0320_), .B(_0245_), .Y(_0346_));
 NAND_g NAND_1373_(.A(_0347_), .B(_0346_), .Y(_0348_));
 NAND_g NAND_1374_(.A(_0301_), .B(SW[6]), .Y(keywire1147));
 NAND_g NAND_1375_(.A(_0328_), .B(_0246_), .Y(_0350_));
 NAND_g NAND_1377_(.A(_0351_), .B(_0348_), .Y(_0160_));
 NAND_g NAND_1378_(.A(_0320_), .B(_0246_), .Y(_0352_));
 NAND_g NAND_1380_(.A(_0353_), .B(_0352_), .Y(_0354_));
 NAND_g NAND_1382_(.A(_0301_), .B(SW[7]), .Y(keywire1148));
 NAND_g NAND_1383_(.A(_0328_), .B(_0247_), .Y(_0357_));
 NAND_g NAND_1385_(.A(_0358_), .B(_0354_), .Y(_0161_));
 NAND_g NAND_1386_(.A(_0301_), .B(SW[8]), .Y(keywire1151));
 NAND_g NAND_1387_(.A(_0321_), .B(T3y[5]), .Y(_0360_));
 NAND_g NAND_1389_(.A(_0361_), .B(_0328_), .Y(_0362_));
 NAND_g NAND_1391_(.A(_0363_), .B(_0360_), .Y(_0162_));
 NAND_g NAND_1392_(.A(_0328_), .B(_0250_), .Y(_0364_));
 NAND_g NAND_1393_(.A(_0320_), .B(_0249_), .Y(_0365_));
 NAND_g NAND_1395_(.A(_0366_), .B(_0365_), .Y(_0367_));
 NAND_g NAND_1396_(.A(_0367_), .B(_0364_), .Y(_0163_));
 NAND_g NAND_1397_(.A(_0301_), .B(SW[0]), .Y(keywire1139));
 NAND_g NAND_1398_(.A(T3plot), .B(T3colourcircle[0]), .Y(_0369_));
 NAND_g NAND_1399_(.A(_0369_), .B(_0368_), .Y(_0164_));
 NAND_g NAND_1400_(.A(_0301_), .B(SW[1]), .Y(keywire1140));
 NAND_g NAND_1401_(.A(T3plot), .B(T3colourcircle[1]), .Y(_0371_));
 NAND_g NAND_1402_(.A(_0371_), .B(_0370_), .Y(_0165_));
 NAND_g NAND_1403_(.A(_0301_), .B(SW[2]), .Y(keywire1141));
 NAND_g NAND_1404_(.A(T3plot), .B(T3colourcircle[2]), .Y(_0373_));
 NAND_g NAND_1405_(.A(_0373_), .B(_0372_), .Y(_0166_));
 NAND_g NAND_1406_(.A(_0303_), .B(_0296_), .Y(_0374_));
 NAND_g NAND_1408_(.A(_0375_), .B(_0253_), .Y(_0376_));
 NAND_g NAND_1410_(.A(1'h1), .B(T3y[0]), .Y(_0378_));
 NAND_g NAND_1412_(.A(_0379_), .B(_0376_), .Y(_0380_));
 NAND_g NAND_1414_(.A(_0264_), .B(_0259_), .Y(_0382_));
 NAND_g NAND_1416_(.A(_0230_), .B(T3x[0]), .Y(_0384_));
 NAND_g NAND_1419_(.A(_0239_), .B(T3xp[0]), .Y(_0387_));
 NAND_g NAND_1420_(.A(_0301_), .B(1'h1), .Y(_0388_));
 NAND_g NAND_1421_(.A(_0388_), .B(_0387_), .Y(_0389_));
 NAND_g NAND_1423_(.A(_0390_), .B(_0380_), .Y(_0167_));
 NAND_g NAND_1424_(.A(1'h1), .B(T3y[1]), .Y(_0391_));
 NAND_g NAND_1427_(.A(_0230_), .B(T3y[0]), .Y(_0394_));
 NAND_g NAND_1428_(.A(_0394_), .B(_0393_), .Y(_0395_));
 NAND_g NAND_1430_(.A(_0396_), .B(_0374_), .Y(_0397_));
 NAND_g NAND_1431_(.A(_0239_), .B(T3xp[1]), .Y(_0398_));
 NAND_g NAND_1432_(.A(_0301_), .B(1'h1), .Y(_0399_));
 NAND_g NAND_1434_(.A(1'h1), .B(T3x[1]), .Y(_0401_));
 NAND_g NAND_1437_(.A(_0403_), .B(_0384_), .Y(_0404_));
 NAND_g NAND_1439_(.A(_0405_), .B(_0305_), .Y(_0406_));
 NAND_g NAND_1441_(.A(1'h1), .B(T3x[0]), .Y(_0408_));
 NAND_g NAND_1442_(.A(_0408_), .B(_0403_), .Y(_0409_));
 NAND_g NAND_1443_(.A(_0407_), .B(_0402_), .Y(_0410_));
 NAND_g NAND_1445_(.A(_0411_), .B(_0410_), .Y(_0412_));
 NAND_g NAND_1446_(.A(_0393_), .B(_0378_), .Y(_0413_));
 NAND_g NAND_1447_(.A(_0392_), .B(_0377_), .Y(_0414_));
 NAND_g NAND_1449_(.A(_0415_), .B(_0414_), .Y(_0416_));
 NAND_g NAND_1453_(.A(_0419_), .B(_0417_), .Y(_0168_));
 NAND_g NAND_1454_(.A(1'h1), .B(T3y[2]), .Y(_0420_));
 NAND_g NAND_1457_(.A(_0414_), .B(_0391_), .Y(_0423_));
 NAND_g NAND_1458_(.A(_0423_), .B(_0421_), .Y(_0424_));
 NAND_g NAND_1460_(.A(_0425_), .B(_0252_), .Y(_0426_));
 NAND_g NAND_1461_(.A(_0239_), .B(T3xp[2]), .Y(_0427_));
 NAND_g NAND_1462_(.A(_0301_), .B(1'h1), .Y(_0428_));
 NAND_g NAND_1465_(.A(1'h1), .B(_0214_), .Y(_0431_));
 NAND_g NAND_1466_(.A(_0431_), .B(_0395_), .Y(_0432_));
 NAND_g NAND_1467_(.A(_0432_), .B(_0422_), .Y(_0433_));
 NAND_g NAND_1469_(.A(_0434_), .B(_0374_), .Y(_0435_));
 NAND_g NAND_1470_(.A(1'h1), .B(T3x[2]), .Y(_0436_));
 NAND_g NAND_1474_(.A(_0410_), .B(_0401_), .Y(_0440_));
 NAND_g NAND_1475_(.A(_0440_), .B(_0437_), .Y(_0441_));
 NAND_g NAND_1476_(.A(_0439_), .B(_0438_), .Y(_0442_));
 NAND_g NAND_1478_(.A(_0443_), .B(_0441_), .Y(_0444_));
 NAND_g NAND_1479_(.A(1'h1), .B(_0222_), .Y(_0445_));
 NAND_g NAND_1481_(.A(_0445_), .B(_0404_), .Y(_0447_));
 NAND_g NAND_1482_(.A(_0446_), .B(_0437_), .Y(_0448_));
 NAND_g NAND_1483_(.A(_0447_), .B(_0438_), .Y(_0449_));
 NAND_g NAND_1485_(.A(_0450_), .B(_0448_), .Y(_0451_));
 NAND_g NAND_1488_(.A(_0453_), .B(_0452_), .Y(_0169_));
 NAND_g NAND_1489_(.A(_0239_), .B(T3xp[3]), .Y(_0454_));
 NAND_g NAND_1490_(.A(_0301_), .B(1'h1), .Y(_0455_));
 NAND_g NAND_1492_(.A(_0231_), .B(_0216_), .Y(_0457_));
 NAND_g NAND_1493_(.A(1'h1), .B(T3y[3]), .Y(_0458_));
 NAND_g NAND_1497_(.A(_0461_), .B(_0252_), .Y(_0462_));
 NAND_g NAND_1498_(.A(_0231_), .B(_0224_), .Y(_0463_));
 NAND_g NAND_1499_(.A(1'h1), .B(T3x[3]), .Y(_0464_));
 NAND_g NAND_1501_(.A(1'h1), .B(_0223_), .Y(_0466_));
 NAND_g NAND_1502_(.A(_0466_), .B(_0449_), .Y(_0467_));
 NAND_g NAND_1504_(.A(_0468_), .B(_0305_), .Y(_0469_));
 NAND_g NAND_1505_(.A(1'h1), .B(_0215_), .Y(_0470_));
 NAND_g NAND_1508_(.A(_0472_), .B(_0374_), .Y(_0473_));
 NAND_g NAND_1511_(.A(_0475_), .B(_0260_), .Y(_0476_));
 NAND_g NAND_1515_(.A(_0479_), .B(_0477_), .Y(_0170_));
 NAND_g NAND_1516_(.A(1'h0), .B(T3y[4]), .Y(_0480_));
 NAND_g NAND_1519_(.A(_0460_), .B(_0458_), .Y(_0483_));
 NAND_g NAND_1521_(.A(_0484_), .B(_0481_), .Y(_0485_));
 NAND_g NAND_1523_(.A(_0486_), .B(_0252_), .Y(_0487_));
 NAND_g NAND_1524_(.A(1'h0), .B(T3x[4]), .Y(_0488_));
 NAND_g NAND_1527_(.A(_0474_), .B(_0464_), .Y(_0491_));
 NAND_g NAND_1530_(.A(_0492_), .B(_0489_), .Y(_0494_));
 NAND_g NAND_1531_(.A(_0494_), .B(_0260_), .Y(_0495_));
 NAND_g NAND_1533_(.A(_0239_), .B(T3xp[4]), .Y(_0497_));
 NAND_g NAND_1534_(.A(_0301_), .B(1'h0), .Y(_0498_));
 NAND_g NAND_1535_(.A(_0498_), .B(_0497_), .Y(_0499_));
 NAND_g NAND_1538_(.A(_0231_), .B(T3x[3]), .Y(_0502_));
 NAND_g NAND_1539_(.A(1'h1), .B(_0224_), .Y(_0503_));
 NAND_g NAND_1540_(.A(_0502_), .B(_0467_), .Y(_0504_));
 NAND_g NAND_1541_(.A(_0504_), .B(_0503_), .Y(_0505_));
 NAND_g NAND_1543_(.A(_0506_), .B(_0489_), .Y(_0507_));
 NAND_g NAND_1544_(.A(_0505_), .B(_0490_), .Y(_0508_));
 NAND_g NAND_1546_(.A(_0509_), .B(_0507_), .Y(_0510_));
 NAND_g NAND_1547_(.A(_0231_), .B(T3y[3]), .Y(_0511_));
 NAND_g NAND_1548_(.A(1'h1), .B(_0216_), .Y(_0512_));
 NAND_g NAND_1549_(.A(_0512_), .B(_0471_), .Y(_0513_));
 NAND_g NAND_1551_(.A(_0514_), .B(_0482_), .Y(_0515_));
 NAND_g NAND_1553_(.A(_0516_), .B(_0374_), .Y(_0517_));
 NAND_g NAND_1555_(.A(_0518_), .B(_0501_), .Y(_0171_));
 NAND_g NAND_1556_(.A(_0232_), .B(_0226_), .Y(_0519_));
 NAND_g NAND_1557_(.A(1'h0), .B(T3x[5]), .Y(_0520_));
 NAND_g NAND_1559_(.A(1'h0), .B(_0225_), .Y(_0522_));
 NAND_g NAND_1560_(.A(_0522_), .B(_0508_), .Y(_0523_));
 NAND_g NAND_1562_(.A(_0232_), .B(_0218_), .Y(_0525_));
 NAND_g NAND_1563_(.A(1'h0), .B(T3y[5]), .Y(_0526_));
 NAND_g NAND_1567_(.A(_0529_), .B(_0252_), .Y(_0530_));
 NAND_g NAND_1568_(.A(_0239_), .B(T3xp[5]), .Y(_0531_));
 NAND_g NAND_1569_(.A(_0301_), .B(1'h0), .Y(_0532_));
 NAND_g NAND_1571_(.A(1'h0), .B(_0217_), .Y(_0534_));
 NAND_g NAND_1574_(.A(_0536_), .B(_0374_), .Y(_0537_));
 NAND_g NAND_1577_(.A(_0539_), .B(_0260_), .Y(_0540_));
 NAND_g NAND_1579_(.A(_0541_), .B(_0305_), .Y(_0542_));
 NAND_g NAND_1582_(.A(_0544_), .B(_0538_), .Y(_0172_));
 NAND_g NAND_1583_(.A(1'h1), .B(T3x[6]), .Y(_0545_));
 NAND_g NAND_1586_(.A(_0524_), .B(_0520_), .Y(_0548_));
 NAND_g NAND_1588_(.A(_0549_), .B(_0546_), .Y(_0550_));
 NAND_g NAND_1590_(.A(_0551_), .B(_0260_), .Y(_0552_));
 NAND_g NAND_1591_(.A(_0301_), .B(1'h1), .Y(_0553_));
 NAND_g NAND_1592_(.A(_0239_), .B(T3xp[6]), .Y(_0554_));
 NAND_g NAND_1594_(.A(1'h1), .B(T3y[6]), .Y(_0556_));
 NAND_g NAND_1597_(.A(_0528_), .B(_0526_), .Y(_0559_));
 NAND_g NAND_1599_(.A(_0560_), .B(_0557_), .Y(_0561_));
 NAND_g NAND_1601_(.A(_0562_), .B(_0252_), .Y(_0563_));
 NAND_g NAND_1604_(.A(1'h0), .B(_0218_), .Y(_0566_));
 NAND_g NAND_1605_(.A(_0232_), .B(T3y[5]), .Y(_0567_));
 NAND_g NAND_1606_(.A(_0566_), .B(_0535_), .Y(_0568_));
 NAND_g NAND_1608_(.A(_0569_), .B(_0558_), .Y(_0570_));
 NAND_g NAND_1610_(.A(_0571_), .B(_0374_), .Y(_0572_));
 NAND_g NAND_1611_(.A(1'h0), .B(_0226_), .Y(_0573_));
 NAND_g NAND_1612_(.A(_0232_), .B(T3x[5]), .Y(_0574_));
 NAND_g NAND_1613_(.A(_0574_), .B(_0523_), .Y(_0575_));
 NAND_g NAND_1615_(.A(_0575_), .B(_0573_), .Y(_0577_));
 NAND_g NAND_1616_(.A(_0577_), .B(_0547_), .Y(_0578_));
 NAND_g NAND_1617_(.A(_0576_), .B(_0546_), .Y(_0579_));
 NAND_g NAND_1619_(.A(_0580_), .B(_0578_), .Y(_0581_));
 NAND_g NAND_1621_(.A(_0582_), .B(_0565_), .Y(_0173_));
 NAND_g NAND_1624_(.A(_0584_), .B(_0252_), .Y(_0585_));
 NAND_g NAND_1625_(.A(_0239_), .B(T3xp[7]), .Y(_0586_));
 NAND_g NAND_1626_(.A(_0301_), .B(1'h0), .Y(_0587_));
 NAND_g NAND_1631_(.A(_0591_), .B(_0260_), .Y(_0592_));
 NAND_g NAND_1632_(.A(1'h1), .B(_0227_), .Y(_0593_));
 NAND_g NAND_1633_(.A(_0593_), .B(_0578_), .Y(_0594_));
 NAND_g NAND_1635_(.A(_0595_), .B(_0305_), .Y(_0596_));
 NAND_g NAND_1636_(.A(1'h1), .B(_0219_), .Y(_0597_));
 NAND_g NAND_1637_(.A(_0597_), .B(_0570_), .Y(_0598_));
 NAND_g NAND_1639_(.A(_0599_), .B(_0374_), .Y(_0600_));
 NAND_g NAND_1643_(.A(_0603_), .B(_0601_), .Y(_0174_));
 NAND_g NAND_1646_(.A(_0326_), .B(_0301_), .Y(_0605_));
 NAND_g NAND_1650_(.A(_0608_), .B(_0605_), .Y(_0176_));
 NAND_g NAND_1651_(.A(T3x[0]), .B(T3y[0]), .Y(_0609_));
 NAND_g NAND_1657_(.A(_0614_), .B(_0319_), .Y(_0615_));
 NAND_g NAND_1658_(.A(_0612_), .B(_0318_), .Y(_0616_));
 NAND_g NAND_1659_(.A(_0616_), .B(_0615_), .Y(_0617_));
 NAND_g NAND_1661_(.A(_0617_), .B(_0607_), .Y(_0619_));
 NAND_g NAND_1663_(.A(_0620_), .B(_0618_), .Y(_0621_));
 NAND_g NAND_1664_(.A(_0238_), .B(T3d[2]), .Y(_0622_));
 NAND_g NAND_1667_(.A(_0624_), .B(_0619_), .Y(_0177_));
 NAND_g NAND_1669_(.A(_0612_), .B(T3d[1]), .Y(_0626_));
 NAND_g NAND_1672_(.A(_0628_), .B(_0214_), .Y(_0629_));
 NAND_g NAND_1674_(.A(_0630_), .B(_0609_), .Y(_0631_));
 NAND_g NAND_1676_(.A(_0632_), .B(T3d[3]), .Y(_0633_));
 NAND_g NAND_1678_(.A(_0634_), .B(_0611_), .Y(_0635_));
 NAND_g NAND_1680_(.A(_0636_), .B(_0626_), .Y(_0637_));
 NAND_g NAND_1681_(.A(_0634_), .B(_0625_), .Y(_0638_));
 NAND_g NAND_1682_(.A(_0614_), .B(_0220_), .Y(_0639_));
 NAND_g NAND_1683_(.A(_0628_), .B(T3d[3]), .Y(_0640_));
 NAND_g NAND_1685_(.A(_0641_), .B(_0613_), .Y(_0642_));
 NAND_g NAND_1692_(.A(_0648_), .B(_0637_), .Y(_0649_));
 NAND_g NAND_1693_(.A(_0649_), .B(_0647_), .Y(_0650_));
 NAND_g NAND_1699_(.A(_0655_), .B(_0650_), .Y(_0178_));
 NAND_g NAND_1700_(.A(_0635_), .B(_0633_), .Y(_0656_));
 NAND_g NAND_1701_(.A(_0631_), .B(_0629_), .Y(_0657_));
 NAND_g NAND_1704_(.A(_0659_), .B(_0215_), .Y(_0660_));
 NAND_g NAND_1706_(.A(_0661_), .B(_0657_), .Y(_0662_));
 NAND_g NAND_1708_(.A(_0663_), .B(T3d[4]), .Y(_0664_));
 NAND_g NAND_1710_(.A(_0665_), .B(_0656_), .Y(_0666_));
 NAND_g NAND_1714_(.A(_0669_), .B(_0318_), .Y(_0670_));
 NAND_g NAND_1715_(.A(_0642_), .B(_0640_), .Y(_0671_));
 NAND_g NAND_1716_(.A(_0659_), .B(T3d[4]), .Y(_0672_));
 NAND_g NAND_1718_(.A(_0673_), .B(_0671_), .Y(_0674_));
 NAND_g NAND_1724_(.A(_0679_), .B(_0677_), .Y(_0680_));
 NAND_g NAND_1725_(.A(_0680_), .B(_0670_), .Y(_0681_));
 NAND_g NAND_1726_(.A(_0681_), .B(_0295_), .Y(_0682_));
 NAND_g NAND_1727_(.A(_0238_), .B(T3d[4]), .Y(_0683_));
 NAND_g NAND_1731_(.A(_0686_), .B(_0682_), .Y(_0179_));
 NAND_g NAND_1732_(.A(_0666_), .B(_0664_), .Y(_0687_));
 NAND_g NAND_1733_(.A(_0662_), .B(_0660_), .Y(_0688_));
 NAND_g NAND_1737_(.A(_0690_), .B(_0216_), .Y(_0692_));
 NAND_g NAND_1738_(.A(_0691_), .B(T3y[3]), .Y(_0693_));
 NAND_g NAND_1741_(.A(_0695_), .B(T3d[5]), .Y(_0696_));
 NAND_g NAND_1743_(.A(_0697_), .B(_0687_), .Y(_0698_));
 NAND_g NAND_1747_(.A(_0701_), .B(_0318_), .Y(_0702_));
 NAND_g NAND_1748_(.A(_0674_), .B(_0672_), .Y(_0703_));
 NAND_g NAND_1749_(.A(_0690_), .B(T3d[5]), .Y(_0704_));
 NAND_g NAND_1751_(.A(_0705_), .B(_0703_), .Y(_0706_));
 NAND_g NAND_1755_(.A(_0709_), .B(_0319_), .Y(_0710_));
 NAND_g NAND_1756_(.A(_0710_), .B(_0702_), .Y(_0711_));
 NAND_g NAND_1757_(.A(_0711_), .B(_0295_), .Y(_0712_));
 NAND_g NAND_1758_(.A(_0238_), .B(T3d[5]), .Y(_0713_));
 NAND_g NAND_1762_(.A(_0716_), .B(_0712_), .Y(_0180_));
 NAND_g NAND_1763_(.A(_0698_), .B(_0696_), .Y(_0717_));
 NAND_g NAND_1766_(.A(_0719_), .B(_0217_), .Y(_0720_));
 NAND_g NAND_1768_(.A(_0693_), .B(_0688_), .Y(_0722_));
 NAND_g NAND_1769_(.A(_0722_), .B(_0692_), .Y(_0723_));
 NAND_g NAND_1770_(.A(_0723_), .B(_0721_), .Y(_0724_));
 NAND_g NAND_1772_(.A(_0725_), .B(T3d[6]), .Y(_0726_));
 NAND_g NAND_1774_(.A(_0727_), .B(_0717_), .Y(_0728_));
 NAND_g NAND_1778_(.A(_0731_), .B(_0318_), .Y(_0732_));
 NAND_g NAND_1779_(.A(_0706_), .B(_0704_), .Y(_0733_));
 NAND_g NAND_1780_(.A(_0719_), .B(T3d[6]), .Y(_0734_));
 NAND_g NAND_1782_(.A(_0735_), .B(_0733_), .Y(_0736_));
 NAND_g NAND_1788_(.A(_0741_), .B(_0739_), .Y(_0742_));
 NAND_g NAND_1789_(.A(_0742_), .B(_0732_), .Y(_0743_));
 NAND_g NAND_1790_(.A(_0743_), .B(_0295_), .Y(_0744_));
 NAND_g NAND_1791_(.A(_0238_), .B(T3d[6]), .Y(_0745_));
 NAND_g NAND_1795_(.A(_0748_), .B(_0744_), .Y(_0181_));
 NAND_g NAND_1796_(.A(_0728_), .B(_0726_), .Y(_0749_));
 NAND_g NAND_1797_(.A(_0724_), .B(_0720_), .Y(_0750_));
 NAND_g NAND_1801_(.A(_0752_), .B(_0218_), .Y(_0754_));
 NAND_g NAND_1802_(.A(_0753_), .B(T3y[5]), .Y(_0755_));
 NAND_g NAND_1805_(.A(_0757_), .B(T3d[7]), .Y(_0758_));
 NAND_g NAND_1807_(.A(_0759_), .B(_0749_), .Y(_0760_));
 NAND_g NAND_1811_(.A(_0763_), .B(_0318_), .Y(_0764_));
 NAND_g NAND_1812_(.A(_0736_), .B(_0734_), .Y(_0765_));
 NAND_g NAND_1813_(.A(_0752_), .B(T3d[7]), .Y(_0766_));
 NAND_g NAND_1815_(.A(_0767_), .B(_0765_), .Y(_0768_));
 NAND_g NAND_1818_(.A(_0769_), .B(_0738_), .Y(_0771_));
 NAND_g NAND_1820_(.A(_0772_), .B(_0771_), .Y(_0773_));
 NAND_g NAND_1821_(.A(_0773_), .B(_0764_), .Y(_0774_));
 NAND_g NAND_1822_(.A(_0774_), .B(_0295_), .Y(_0775_));
 NAND_g NAND_1823_(.A(_0238_), .B(T3d[7]), .Y(_0776_));
 NAND_g NAND_1825_(.A(_0777_), .B(_0775_), .Y(_0182_));
 NAND_g NAND_1826_(.A(_0760_), .B(_0758_), .Y(_0778_));
 NAND_g NAND_1827_(.A(_0755_), .B(_0750_), .Y(_0779_));
 NAND_g NAND_1836_(.A(_0787_), .B(_0318_), .Y(_0788_));
 NAND_g NAND_1837_(.A(_0768_), .B(_0766_), .Y(_0789_));
 NAND_g NAND_1840_(.A(_0791_), .B(_0319_), .Y(_0792_));
 NAND_g NAND_1841_(.A(_0792_), .B(_0788_), .Y(_0793_));
 NAND_g NAND_1842_(.A(_0793_), .B(_0295_), .Y(_0794_));
 NAND_g NAND_1843_(.A(_0238_), .B(T3d[8]), .Y(_0795_));
 NAND_g NAND_1845_(.A(_0796_), .B(_0794_), .Y(_0183_));
 NAND_g NAND_1846_(.A(_0238_), .B(T3x[0]), .Y(_0797_));
 NAND_g NAND_1847_(.A(_0295_), .B(_0221_), .Y(_0798_));
 NAND_g NAND_1848_(.A(_0798_), .B(_0797_), .Y(_0184_));
 NAND_g NAND_1849_(.A(_0238_), .B(T3x[1]), .Y(_0799_));
 NAND_g NAND_1850_(.A(_0628_), .B(_0295_), .Y(_0800_));
 NAND_g NAND_1851_(.A(_0800_), .B(_0799_), .Y(_0185_));
 NAND_g NAND_1852_(.A(_0238_), .B(T3x[2]), .Y(_0801_));
 NAND_g NAND_1853_(.A(_0659_), .B(_0295_), .Y(_0802_));
 NAND_g NAND_1854_(.A(_0802_), .B(_0801_), .Y(_0186_));
 NAND_g NAND_1855_(.A(_0238_), .B(T3x[3]), .Y(_0803_));
 NAND_g NAND_1856_(.A(_0690_), .B(_0295_), .Y(_0804_));
 NAND_g NAND_1857_(.A(_0804_), .B(_0803_), .Y(_0187_));
 NAND_g NAND_1858_(.A(_0238_), .B(T3x[4]), .Y(_0805_));
 NAND_g NAND_1859_(.A(_0719_), .B(_0295_), .Y(_0806_));
 NAND_g NAND_1860_(.A(_0806_), .B(_0805_), .Y(_0188_));
 NAND_g NAND_1861_(.A(_0238_), .B(T3x[5]), .Y(_0807_));
 NAND_g NAND_1862_(.A(_0752_), .B(_0295_), .Y(_0808_));
 NAND_g NAND_1863_(.A(_0808_), .B(_0807_), .Y(_0189_));
 NAND_g NAND_1864_(.A(_0238_), .B(T3x[6]), .Y(_0809_));
 NAND_g NAND_1865_(.A(_0782_), .B(_0295_), .Y(_0810_));
 NAND_g NAND_1866_(.A(_0810_), .B(_0809_), .Y(_0190_));
 NAND_g NAND_1867_(.A(_0781_), .B(_0297_), .Y(_0811_));
 NAND_g NAND_1868_(.A(_0781_), .B(_0237_), .Y(_0812_));
 NAND_g NAND_1870_(.A(_0813_), .B(_0812_), .Y(_0814_));
 NAND_g NAND_1871_(.A(_0814_), .B(_0811_), .Y(_0191_));
 NAND_g NAND_1873_(.A(_0233_), .B(T3y[0]), .Y(_0816_));
 NAND_g NAND_1885_(.A(_0827_), .B(_0820_), .Y(_0192_));
 NAND_g NAND_1887_(.A(_0336_), .B(1'h1), .Y(_0829_));
 NAND_g NAND_1889_(.A(_0830_), .B(_0828_), .Y(_0831_));
 NAND_g NAND_1891_(.A(_0832_), .B(_0301_), .Y(_0833_));
 NAND_g NAND_1892_(.A(_0239_), .B(T3yp[1]), .Y(_0834_));
 NAND_g NAND_1893_(.A(1'h1), .B(T3y[1]), .Y(_0835_));
 NAND_g NAND_1896_(.A(_0836_), .B(_0815_), .Y(_0838_));
 NAND_g NAND_1898_(.A(_0839_), .B(_0381_), .Y(_0840_));
 NAND_g NAND_1899_(.A(1'h1), .B(T3x[1]), .Y(_0841_));
 NAND_g NAND_1902_(.A(_0842_), .B(_0821_), .Y(_0844_));
 NAND_g NAND_1904_(.A(_0845_), .B(_0265_), .Y(_0846_));
 NAND_g NAND_1905_(.A(_0837_), .B(_0816_), .Y(_0847_));
 NAND_g NAND_1907_(.A(_0848_), .B(_0262_), .Y(_0849_));
 NAND_g NAND_1908_(.A(_0296_), .B(_0254_), .Y(_0850_));
 NAND_g NAND_1909_(.A(_0233_), .B(T3x[0]), .Y(_0851_));
 NAND_g NAND_1910_(.A(_0851_), .B(_0843_), .Y(_0852_));
 NAND_g NAND_1912_(.A(_0853_), .B(_0850_), .Y(_0854_));
 NAND_g NAND_1917_(.A(_0858_), .B(_0833_), .Y(_0193_));
 NAND_g NAND_1918_(.A(_0831_), .B(_0829_), .Y(_0859_));
 NAND_g NAND_1919_(.A(_0342_), .B(1'h0), .Y(_0860_));
 NAND_g NAND_1921_(.A(_0861_), .B(_0859_), .Y(_0862_));
 NAND_g NAND_1923_(.A(_0863_), .B(_0301_), .Y(_0864_));
 NAND_g NAND_1924_(.A(1'h0), .B(T3x[2]), .Y(_0865_));
 NAND_g NAND_1928_(.A(_0844_), .B(_0841_), .Y(_0869_));
 NAND_g NAND_1929_(.A(_0869_), .B(_0866_), .Y(_0870_));
 NAND_g NAND_1930_(.A(_0868_), .B(_0867_), .Y(_0871_));
 NAND_g NAND_1932_(.A(_0872_), .B(_0870_), .Y(_0873_));
 NAND_g NAND_1933_(.A(_0239_), .B(T3yp[2]), .Y(_0874_));
 NAND_g NAND_1935_(.A(1'h1), .B(_0222_), .Y(_0876_));
 NAND_g NAND_1936_(.A(_0876_), .B(_0852_), .Y(_0877_));
 NAND_g NAND_1937_(.A(_0877_), .B(_0867_), .Y(_0878_));
 NAND_g NAND_1939_(.A(_0879_), .B(_0850_), .Y(_0880_));
 NAND_g NAND_1940_(.A(1'h0), .B(T3y[2]), .Y(_0881_));
 NAND_g NAND_1943_(.A(1'h1), .B(_0214_), .Y(_0884_));
 NAND_g NAND_1944_(.A(_0884_), .B(_0847_), .Y(_0885_));
 NAND_g NAND_1945_(.A(_0885_), .B(_0883_), .Y(_0886_));
 NAND_g NAND_1947_(.A(_0887_), .B(_0262_), .Y(_0888_));
 NAND_g NAND_1949_(.A(_0838_), .B(_0835_), .Y(_0890_));
 NAND_g NAND_1950_(.A(_0889_), .B(_0883_), .Y(_0891_));
 NAND_g NAND_1951_(.A(_0890_), .B(_0882_), .Y(_0892_));
 NAND_g NAND_1953_(.A(_0893_), .B(_0891_), .Y(_0894_));
 NAND_g NAND_1957_(.A(_0897_), .B(_0864_), .Y(_0194_));
 NAND_g NAND_1958_(.A(_0862_), .B(_0860_), .Y(_0898_));
 NAND_g NAND_1963_(.A(_0902_), .B(_0301_), .Y(_0903_));
 NAND_g NAND_1964_(.A(_0234_), .B(_0224_), .Y(_0904_));
 NAND_g NAND_1965_(.A(1'h1), .B(T3x[3]), .Y(_0905_));
 NAND_g NAND_1967_(.A(1'h0), .B(_0223_), .Y(_0907_));
 NAND_g NAND_1968_(.A(_0907_), .B(_0878_), .Y(_0908_));
 NAND_g NAND_1970_(.A(_0908_), .B(_0850_), .Y(_0910_));
 NAND_g NAND_1973_(.A(_0911_), .B(_0265_), .Y(_0913_));
 NAND_g NAND_1974_(.A(_0913_), .B(_0910_), .Y(_0914_));
 NAND_g NAND_1975_(.A(_0914_), .B(_0906_), .Y(_0915_));
 NAND_g NAND_1976_(.A(_0239_), .B(T3yp[3]), .Y(_0916_));
 NAND_g NAND_1977_(.A(_0234_), .B(_0216_), .Y(_0917_));
 NAND_g NAND_1978_(.A(1'h1), .B(T3y[3]), .Y(_0918_));
 NAND_g NAND_1980_(.A(1'h0), .B(_0215_), .Y(_0920_));
 NAND_g NAND_1981_(.A(_0920_), .B(_0886_), .Y(_0921_));
 NAND_g NAND_1983_(.A(_0922_), .B(_0262_), .Y(_0923_));
 NAND_g NAND_1986_(.A(_0925_), .B(_0381_), .Y(_0926_));
 NAND_g NAND_1989_(.A(_0909_), .B(_0850_), .Y(_0929_));
 NAND_g NAND_1990_(.A(_0912_), .B(_0265_), .Y(_0930_));
 NAND_g NAND_1993_(.A(_0921_), .B(_0262_), .Y(_0933_));
 NAND_g NAND_1994_(.A(_0924_), .B(_0381_), .Y(_0934_));
 NAND_g NAND_1995_(.A(_0934_), .B(_0933_), .Y(_0935_));
 NAND_g NAND_1996_(.A(_0935_), .B(_0919_), .Y(_0936_));
 NAND_g NAND_2001_(.A(_0940_), .B(_0903_), .Y(_0195_));
 NAND_g NAND_2002_(.A(_0355_), .B(1'h1), .Y(_0941_));
 NAND_g NAND_2006_(.A(_0944_), .B(_0942_), .Y(_0945_));
 NAND_g NAND_2008_(.A(_0946_), .B(_0301_), .Y(_0947_));
 NAND_g NAND_2009_(.A(1'h1), .B(T3x[4]), .Y(_0948_));
 NAND_g NAND_2012_(.A(_0234_), .B(T3x[3]), .Y(_0951_));
 NAND_g NAND_2013_(.A(1'h1), .B(_0224_), .Y(_0952_));
 NAND_g NAND_2014_(.A(_0951_), .B(_0908_), .Y(_0953_));
 NAND_g NAND_2015_(.A(_0953_), .B(_0952_), .Y(_0954_));
 NAND_g NAND_2016_(.A(_0954_), .B(_0950_), .Y(_0955_));
 NAND_g NAND_2018_(.A(_0956_), .B(_0850_), .Y(_0957_));
 NAND_g NAND_2019_(.A(1'h1), .B(T3y[4]), .Y(_0958_));
 NAND_g NAND_2022_(.A(_0234_), .B(T3y[3]), .Y(_0961_));
 NAND_g NAND_2023_(.A(1'h1), .B(_0216_), .Y(_0962_));
 NAND_g NAND_2024_(.A(_0961_), .B(_0921_), .Y(_0963_));
 NAND_g NAND_2025_(.A(_0963_), .B(_0962_), .Y(_0964_));
 NAND_g NAND_2026_(.A(_0964_), .B(_0960_), .Y(_0965_));
 NAND_g NAND_2028_(.A(_0966_), .B(_0262_), .Y(_0967_));
 NAND_g NAND_2030_(.A(_0911_), .B(_0905_), .Y(_0969_));
 NAND_g NAND_2033_(.A(_0970_), .B(_0949_), .Y(_0972_));
 NAND_g NAND_2034_(.A(_0972_), .B(_0265_), .Y(_0973_));
 NAND_g NAND_2036_(.A(_0239_), .B(T3yp[4]), .Y(_0975_));
 NAND_g NAND_2037_(.A(_0924_), .B(_0918_), .Y(_0976_));
 NAND_g NAND_2040_(.A(_0977_), .B(_0959_), .Y(_0979_));
 NAND_g NAND_2042_(.A(_0980_), .B(_0979_), .Y(_0981_));
 NAND_g NAND_2043_(.A(_0981_), .B(_0975_), .Y(_0982_));
 NAND_g NAND_2046_(.A(_0984_), .B(_0947_), .Y(_0196_));
 NAND_g NAND_2047_(.A(_0945_), .B(_0941_), .Y(_0985_));
 NAND_g NAND_2049_(.A(_0359_), .B(_0235_), .Y(_0987_));
 NAND_g NAND_2052_(.A(_0989_), .B(_0301_), .Y(_0990_));
 NAND_g NAND_2053_(.A(_0235_), .B(_0226_), .Y(_0991_));
 NAND_g NAND_2054_(.A(1'h1), .B(T3x[5]), .Y(_0992_));
 NAND_g NAND_2058_(.A(_0995_), .B(_0265_), .Y(_0996_));
 NAND_g NAND_2059_(.A(_0239_), .B(T3yp[5]), .Y(_0997_));
 NAND_g NAND_2060_(.A(_0235_), .B(T3y[5]), .Y(_0998_));
 NAND_g NAND_2061_(.A(1'h1), .B(_0218_), .Y(_0999_));
 NAND_g NAND_2062_(.A(_0235_), .B(_0218_), .Y(_1000_));
 NAND_g NAND_2063_(.A(1'h1), .B(T3y[5]), .Y(_1001_));
 NAND_g NAND_2067_(.A(_1004_), .B(_0381_), .Y(_1005_));
 NAND_g NAND_2070_(.A(1'h1), .B(_0225_), .Y(_1008_));
 NAND_g NAND_2073_(.A(_1010_), .B(_0850_), .Y(_1011_));
 NAND_g NAND_2074_(.A(1'h1), .B(_0217_), .Y(_1012_));
 NAND_g NAND_2075_(.A(_1012_), .B(_0965_), .Y(_1013_));
 NAND_g NAND_2077_(.A(_1014_), .B(_0262_), .Y(_1015_));
 NAND_g NAND_2080_(.A(_1017_), .B(_0990_), .Y(_0197_));
 NAND_g NAND_2084_(.A(_1020_), .B(_0301_), .Y(_1021_));
 NAND_g NAND_2085_(.A(_1003_), .B(_1001_), .Y(_1022_));
 NAND_g NAND_2089_(.A(_1025_), .B(_0381_), .Y(_1026_));
 NAND_g NAND_2090_(.A(_0239_), .B(T3yp[6]), .Y(_1027_));
 NAND_g NAND_2093_(.A(_0994_), .B(_0992_), .Y(_1030_));
 NAND_g NAND_2095_(.A(_1031_), .B(_1029_), .Y(_1032_));
 NAND_g NAND_2097_(.A(_1032_), .B(_0265_), .Y(_1034_));
 NAND_g NAND_2099_(.A(_1013_), .B(_0998_), .Y(_1036_));
 NAND_g NAND_2102_(.A(_0199_), .B(_0262_), .Y(_0200_));
 NAND_g NAND_2103_(.A(1'h1), .B(_0226_), .Y(_0201_));
 NAND_g NAND_2104_(.A(_0235_), .B(T3x[5]), .Y(_0202_));
 NAND_g NAND_2105_(.A(_0201_), .B(_1009_), .Y(_0203_));
 NAND_g NAND_2112_(.A(_0209_), .B(_1021_), .Y(_0198_));
 AND_g AND_1101_(.A(T2x[0]), .B(T2x[1]), .Y(keywire1157));
 AND_g AND_1102_(.A(_0116_), .B(T2x[2]), .Y(keywire1161));
 AND_g AND_1103_(.A(_0117_), .B(T2x[3]), .Y(keywire1164));
 AND_g AND_1104_(.A(_0118_), .B(T2x[4]), .Y(keywire1167));
 AND_g AND_1106_(.A(_0120_), .B(T2x[7]), .Y(_0121_));
 AND_g AND_1107_(.A(_0121_), .B(_0119_), .Y(_0122_));
 AND_g AND_1109_(.A(T2y[0]), .B(T2y[1]), .Y(_0124_));
 AND_g AND_1110_(.A(_0124_), .B(T2y[2]), .Y(_0125_));
 AND_g AND_1111_(.A(T2y[5]), .B(T2y[6]), .Y(_0126_));
 AND_g AND_1114_(.A(_0128_), .B(_0125_), .Y(_0129_));
 AND_g AND_1120_(.A(_0125_), .B(T2y[3]), .Y(_0134_));
 AND_g AND_1121_(.A(_0134_), .B(T2y[4]), .Y(_0135_));
 AND_g AND_1122_(.A(_0135_), .B(T2y[5]), .Y(_0136_));
 AND_g AND_1125_(.A(_0138_), .B(T2x[7]), .Y(_0139_));
 AND_g AND_1128_(.A(_0136_), .B(_0133_), .Y(_0142_));
 AND_g AND_1155_(.A(_0119_), .B(T2x[5]), .Y(keywire1170));
 AND_g AND_1159_(.A(_0091_), .B(_0141_), .Y(_0063_));
 AND_g AND_1163_(.A(_0093_), .B(_0089_), .Y(_0061_));
 AND_g AND_1177_(.A(_0102_), .B(_0141_), .Y(_0056_));
 AND_g AND_1178_(.A(_0140_), .B(KEY_N[3]), .Y(keywire1138));
 AND_g AND_1180_(.A(_0104_), .B(_0103_), .Y(_0105_));
 AND_g AND_1184_(.A(_0107_), .B(_0103_), .Y(_0108_));
 AND_g AND_1188_(.A(_0110_), .B(_0103_), .Y(_0111_));
 AND_g AND_1254_(.A(_0236_), .B(_0211_), .Y(_0237_));
 AND_g AND_1256_(.A(_0238_), .B(T3state[3]), .Y(_0239_));
 AND_g AND_1258_(.A(_0240_), .B(T2Done), .Y(_0241_));
 AND_g AND_1264_(.A(_0246_), .B(_0217_), .Y(_0247_));
 AND_g AND_1268_(.A(T3state[2]), .B(_0210_), .Y(_0251_));
 AND_g AND_1269_(.A(_0251_), .B(T3state[0]), .Y(_0252_));
 AND_g AND_1278_(.A(_0259_), .B(T3state[0]), .Y(_0260_));
 AND_g AND_1281_(.A(_0212_), .B(T3state[1]), .Y(_0263_));
 AND_g AND_1283_(.A(_0264_), .B(_0251_), .Y(_0265_));
 AND_g AND_1287_(.A(_0268_), .B(_0267_), .Y(_0155_));
 AND_g AND_1289_(.A(_0264_), .B(T2Done), .Y(_0270_));
 AND_g AND_1301_(.A(_0280_), .B(_0279_), .Y(_0281_));
 AND_g AND_1307_(.A(_0286_), .B(_0285_), .Y(_0287_));
 AND_g AND_1311_(.A(_0290_), .B(_0289_), .Y(_0291_));
 AND_g AND_1315_(.A(_0237_), .B(T3state[3]), .Y(_0295_));
 AND_g AND_1319_(.A(_0298_), .B(_0297_), .Y(_0299_));
 AND_g AND_1321_(.A(_0259_), .B(_0236_), .Y(_0301_));
 AND_g AND_1328_(.A(_0306_), .B(_0303_), .Y(_0307_));
 AND_g AND_1335_(.A(_0312_), .B(_0311_), .Y(_0313_));
 AND_g AND_1338_(.A(_0315_), .B(_0314_), .Y(_0316_));
 AND_g AND_1342_(.A(_0318_), .B(_0237_), .Y(_0320_));
 AND_g AND_1345_(.A(SW[6]), .B(SW[5]), .Y(keywire1145));
 AND_g AND_1346_(.A(SW[8]), .B(SW[7]), .Y(keywire1149));
 AND_g AND_1348_(.A(_0325_), .B(_0228_), .Y(_0326_));
 AND_g AND_1350_(.A(_0318_), .B(_0295_), .Y(_0328_));
 AND_g AND_1351_(.A(_0328_), .B(_0213_), .Y(_0329_));
 AND_g AND_1360_(.A(_0335_), .B(_0333_), .Y(_0337_));
 AND_g AND_1363_(.A(T3plot), .B(T3y[2]), .Y(_0339_));
 AND_g AND_1365_(.A(_0301_), .B(SW[5]), .Y(keywire1146));
 AND_g AND_1366_(.A(_0341_), .B(_0325_), .Y(_0342_));
 AND_g AND_1369_(.A(_0344_), .B(_0343_), .Y(_0345_));
 AND_g AND_1372_(.A(T3plot), .B(T3y[3]), .Y(_0347_));
 AND_g AND_1376_(.A(_0350_), .B(_0349_), .Y(_0351_));
 AND_g AND_1379_(.A(T3plot), .B(T3y[4]), .Y(_0353_));
 AND_g AND_1381_(.A(_0301_), .B(SW[7]), .Y(keywire1150));
 AND_g AND_1384_(.A(_0357_), .B(_0356_), .Y(_0358_));
 AND_g AND_1390_(.A(_0362_), .B(_0359_), .Y(_0363_));
 AND_g AND_1394_(.A(T3plot), .B(T3y[6]), .Y(_0366_));
 AND_g AND_1409_(.A(1'h1), .B(T3y[0]), .Y(_0377_));
 AND_g AND_1413_(.A(_0264_), .B(_0259_), .Y(_0381_));
 AND_g AND_1433_(.A(_0399_), .B(_0398_), .Y(_0400_));
 AND_g AND_1440_(.A(1'h1), .B(T3x[0]), .Y(_0407_));
 AND_g AND_1444_(.A(_0409_), .B(_0260_), .Y(_0411_));
 AND_g AND_1448_(.A(_0413_), .B(_0252_), .Y(_0415_));
 AND_g AND_1450_(.A(_0412_), .B(_0406_), .Y(_0417_));
 AND_g AND_1451_(.A(_0416_), .B(_0400_), .Y(_0418_));
 AND_g AND_1452_(.A(_0418_), .B(_0397_), .Y(_0419_));
 AND_g AND_1463_(.A(_0428_), .B(_0427_), .Y(_0429_));
 AND_g AND_1464_(.A(_0429_), .B(_0426_), .Y(_0430_));
 AND_g AND_1473_(.A(_0410_), .B(_0401_), .Y(_0439_));
 AND_g AND_1477_(.A(_0442_), .B(_0260_), .Y(_0443_));
 AND_g AND_1480_(.A(_0445_), .B(_0404_), .Y(_0446_));
 AND_g AND_1484_(.A(_0449_), .B(_0305_), .Y(_0450_));
 AND_g AND_1486_(.A(_0451_), .B(_0435_), .Y(_0452_));
 AND_g AND_1487_(.A(_0444_), .B(_0430_), .Y(_0453_));
 AND_g AND_1491_(.A(_0455_), .B(_0454_), .Y(_0456_));
 AND_g AND_1495_(.A(_0424_), .B(_0420_), .Y(_0460_));
 AND_g AND_1506_(.A(_0470_), .B(_0433_), .Y(_0471_));
 AND_g AND_1509_(.A(_0441_), .B(_0436_), .Y(_0474_));
 AND_g AND_1512_(.A(_0473_), .B(_0456_), .Y(_0477_));
 AND_g AND_1513_(.A(_0469_), .B(_0462_), .Y(_0478_));
 AND_g AND_1514_(.A(_0478_), .B(_0476_), .Y(_0479_));
 AND_g AND_1520_(.A(_0483_), .B(_0457_), .Y(_0484_));
 AND_g AND_1528_(.A(_0491_), .B(_0463_), .Y(_0492_));
 AND_g AND_1537_(.A(_0500_), .B(_0487_), .Y(_0501_));
 AND_g AND_1542_(.A(_0504_), .B(_0503_), .Y(_0506_));
 AND_g AND_1545_(.A(_0508_), .B(_0305_), .Y(_0509_));
 AND_g AND_1550_(.A(_0513_), .B(_0511_), .Y(_0514_));
 AND_g AND_1554_(.A(_0517_), .B(_0510_), .Y(_0518_));
 AND_g AND_1561_(.A(_0494_), .B(_0488_), .Y(_0524_));
 AND_g AND_1565_(.A(_0485_), .B(_0480_), .Y(_0528_));
 AND_g AND_1570_(.A(_0532_), .B(_0531_), .Y(_0533_));
 AND_g AND_1572_(.A(_0534_), .B(_0515_), .Y(_0535_));
 AND_g AND_1575_(.A(_0537_), .B(_0530_), .Y(_0538_));
 AND_g AND_1580_(.A(_0542_), .B(_0533_), .Y(_0543_));
 AND_g AND_1581_(.A(_0543_), .B(_0540_), .Y(_0544_));
 AND_g AND_1587_(.A(_0548_), .B(_0519_), .Y(_0549_));
 AND_g AND_1593_(.A(_0554_), .B(_0553_), .Y(_0555_));
 AND_g AND_1598_(.A(_0559_), .B(_0525_), .Y(_0560_));
 AND_g AND_1602_(.A(_0563_), .B(_0555_), .Y(_0564_));
 AND_g AND_1603_(.A(_0564_), .B(_0552_), .Y(_0565_));
 AND_g AND_1607_(.A(_0568_), .B(_0567_), .Y(_0569_));
 AND_g AND_1614_(.A(_0575_), .B(_0573_), .Y(_0576_));
 AND_g AND_1618_(.A(_0579_), .B(_0305_), .Y(_0580_));
 AND_g AND_1620_(.A(_0581_), .B(_0572_), .Y(_0582_));
 AND_g AND_1622_(.A(_0561_), .B(_0556_), .Y(_0583_));
 AND_g AND_1627_(.A(_0587_), .B(_0586_), .Y(_0588_));
 AND_g AND_1629_(.A(_0550_), .B(_0545_), .Y(_0590_));
 AND_g AND_1640_(.A(_0596_), .B(_0588_), .Y(_0601_));
 AND_g AND_1641_(.A(_0592_), .B(_0585_), .Y(_0602_));
 AND_g AND_1642_(.A(_0602_), .B(_0600_), .Y(_0603_));
 AND_g AND_1647_(.A(_0238_), .B(T3d[1]), .Y(_0606_));
 AND_g AND_1648_(.A(_0295_), .B(_0220_), .Y(_0607_));
 AND_g AND_1653_(.A(_0610_), .B(T3d[2]), .Y(_0611_));
 AND_g AND_1655_(.A(_0221_), .B(T3d[2]), .Y(_0613_));
 AND_g AND_1660_(.A(_0616_), .B(_0615_), .Y(_0618_));
 AND_g AND_1662_(.A(_0295_), .B(T3d[1]), .Y(_0620_));
 AND_g AND_1665_(.A(_0622_), .B(_0335_), .Y(_0623_));
 AND_g AND_1666_(.A(_0623_), .B(_0621_), .Y(_0624_));
 AND_g AND_1668_(.A(_0612_), .B(T3d[1]), .Y(_0625_));
 AND_g AND_1670_(.A(T3x[1]), .B(T3x[0]), .Y(_0627_));
 AND_g AND_1687_(.A(_0643_), .B(_0639_), .Y(_0644_));
 AND_g AND_1691_(.A(_0638_), .B(_0318_), .Y(_0648_));
 AND_g AND_1694_(.A(_0238_), .B(T3d[3]), .Y(_0651_));
 AND_g AND_1695_(.A(_0343_), .B(_0335_), .Y(_0652_));
 AND_g AND_1696_(.A(_0342_), .B(SW[4]), .Y(keywire1144));
 AND_g AND_1702_(.A(_0627_), .B(T3x[2]), .Y(_0658_));
 AND_g AND_1712_(.A(_0667_), .B(_0637_), .Y(_0668_));
 AND_g AND_1720_(.A(_0675_), .B(_0644_), .Y(_0676_));
 AND_g AND_1728_(.A(_0652_), .B(_0349_), .Y(_0684_));
 AND_g AND_1730_(.A(_0685_), .B(_0683_), .Y(_0686_));
 AND_g AND_1734_(.A(_0658_), .B(T3x[3]), .Y(_0689_));
 AND_g AND_1745_(.A(_0699_), .B(_0668_), .Y(_0700_));
 AND_g AND_1753_(.A(_0707_), .B(_0676_), .Y(_0708_));
 AND_g AND_1759_(.A(_0684_), .B(_0356_), .Y(_0714_));
 AND_g AND_1761_(.A(_0715_), .B(_0713_), .Y(_0716_));
 AND_g AND_1764_(.A(_0689_), .B(T3x[4]), .Y(_0718_));
 AND_g AND_1776_(.A(_0729_), .B(_0700_), .Y(_0730_));
 AND_g AND_1784_(.A(_0737_), .B(_0708_), .Y(_0738_));
 AND_g AND_1792_(.A(_0714_), .B(_0359_), .Y(_0746_));
 AND_g AND_1794_(.A(_0747_), .B(_0745_), .Y(_0748_));
 AND_g AND_1798_(.A(_0718_), .B(T3x[5]), .Y(_0751_));
 AND_g AND_1809_(.A(_0761_), .B(_0730_), .Y(_0762_));
 AND_g AND_1824_(.A(_0776_), .B(_0746_), .Y(_0777_));
 AND_g AND_1828_(.A(_0779_), .B(_0754_), .Y(_0780_));
 AND_g AND_1829_(.A(_0751_), .B(T3x[6]), .Y(_0781_));
 AND_g AND_1844_(.A(_0795_), .B(_0746_), .Y(_0796_));
 AND_g AND_1869_(.A(T3plot), .B(T3x[7]), .Y(_0813_));
 AND_g AND_1872_(.A(1'h1), .B(T3y[0]), .Y(_0815_));
 AND_g AND_1876_(.A(_0239_), .B(T3yp[0]), .Y(_0819_));
 AND_g AND_1878_(.A(1'h1), .B(T3x[0]), .Y(_0821_));
 AND_g AND_1880_(.A(_0822_), .B(_0376_), .Y(_0823_));
 AND_g AND_1882_(.A(_0605_), .B(1'h1), .Y(_0825_));
 AND_g AND_1886_(.A(_0327_), .B(1'h1), .Y(_0828_));
 AND_g AND_1913_(.A(_0849_), .B(_0834_), .Y(_0855_));
 AND_g AND_1914_(.A(_0854_), .B(_0846_), .Y(_0856_));
 AND_g AND_1915_(.A(_0856_), .B(_0855_), .Y(_0857_));
 AND_g AND_1916_(.A(_0857_), .B(_0840_), .Y(_0858_));
 AND_g AND_1927_(.A(_0844_), .B(_0841_), .Y(_0868_));
 AND_g AND_1931_(.A(_0871_), .B(_0265_), .Y(_0872_));
 AND_g AND_1934_(.A(_0874_), .B(_0873_), .Y(_0875_));
 AND_g AND_1948_(.A(_0838_), .B(_0835_), .Y(_0889_));
 AND_g AND_1952_(.A(_0892_), .B(_0381_), .Y(_0893_));
 AND_g AND_1954_(.A(_0894_), .B(_0888_), .Y(_0895_));
 AND_g AND_1955_(.A(_0895_), .B(_0880_), .Y(_0896_));
 AND_g AND_1956_(.A(_0896_), .B(_0875_), .Y(_0897_));
 AND_g AND_1960_(.A(_0349_), .B(_0234_), .Y(_0900_));
 AND_g AND_1971_(.A(_0870_), .B(_0865_), .Y(_0911_));
 AND_g AND_1984_(.A(_0892_), .B(_0881_), .Y(_0924_));
 AND_g AND_1987_(.A(_0926_), .B(_0923_), .Y(_0927_));
 AND_g AND_1991_(.A(_0930_), .B(_0929_), .Y(_0931_));
 AND_g AND_1998_(.A(_0936_), .B(_0916_), .Y(_0938_));
 AND_g AND_1999_(.A(_0938_), .B(_0915_), .Y(_0939_));
 AND_g AND_2000_(.A(_0939_), .B(_0937_), .Y(_0940_));
 AND_g AND_2029_(.A(_0967_), .B(_0957_), .Y(_0968_));
 AND_g AND_2031_(.A(_0969_), .B(_0904_), .Y(_0970_));
 AND_g AND_2038_(.A(_0976_), .B(_0917_), .Y(_0977_));
 AND_g AND_2045_(.A(_0983_), .B(_0968_), .Y(_0984_));
 AND_g AND_2056_(.A(_0972_), .B(_0948_), .Y(_0994_));
 AND_g AND_2065_(.A(_0979_), .B(_0958_), .Y(_1003_));
 AND_g AND_2068_(.A(_1005_), .B(_0997_), .Y(_1006_));
 AND_g AND_2069_(.A(_1006_), .B(_0996_), .Y(_1007_));
 AND_g AND_2071_(.A(_1008_), .B(_0955_), .Y(_1009_));
 AND_g AND_2078_(.A(_1015_), .B(_1011_), .Y(_1016_));
 AND_g AND_2079_(.A(_1016_), .B(_1007_), .Y(_1017_));
 AND_g AND_2081_(.A(_0987_), .B(_0985_), .Y(_1018_));
 AND_g AND_2086_(.A(_1022_), .B(_1000_), .Y(_1023_));
 AND_g AND_2091_(.A(_1027_), .B(_1026_), .Y(_1028_));
 AND_g AND_2094_(.A(_1030_), .B(_0991_), .Y(_1031_));
 AND_g AND_2100_(.A(_1036_), .B(_0999_), .Y(_1037_));
 AND_g AND_2106_(.A(_0203_), .B(_0202_), .Y(_0204_));
 AND_g AND_2108_(.A(_0205_), .B(_0850_), .Y(_0206_));
 AND_g AND_2110_(.A(_0207_), .B(_0200_), .Y(_0208_));
 AND_g AND_2111_(.A(_0208_), .B(_1028_), .Y(_0209_));
 NOR_g NOR_1105_(.A(T2x[5]), .B(T2x[6]), .Y(keywire1171));
 NOR_g NOR_1113_(.A(_0127_), .B(T2y[3]), .Y(_0128_));
 NOR_g NOR_1117_(.A(_0125_), .B(T2y[3]), .Y(_0131_));
 NOR_g NOR_1118_(.A(_0131_), .B(_0127_), .Y(_0132_));
 NOR_g NOR_1119_(.A(_0132_), .B(_0123_), .Y(_0133_));
 NOR_g NOR_1123_(.A(_0119_), .B(T2x[5]), .Y(keywire1172));
 NOR_g NOR_1129_(.A(_0142_), .B(T2y[6]), .Y(_0143_));
 NOR_g NOR_1130_(.A(_0141_), .B(_0133_), .Y(_0144_));
 NOR_g NOR_1131_(.A(_0144_), .B(_0143_), .Y(_0070_));
 NOR_g NOR_1160_(.A(_0088_), .B(T2x[6]), .Y(keywire1176));
 NOR_g NOR_1161_(.A(_0092_), .B(_0091_), .Y(_0062_));
 NOR_g NOR_1162_(.A(_0137_), .B(T2x[7]), .Y(_0093_));
 NOR_g NOR_1181_(.A(_0103_), .B(T2colour[0]), .Y(_0106_));
 NOR_g NOR_1182_(.A(_0106_), .B(_0105_), .Y(_0072_));
 NOR_g NOR_1185_(.A(_0103_), .B(T2colour[1]), .Y(_0109_));
 NOR_g NOR_1186_(.A(_0109_), .B(_0108_), .Y(_0073_));
 NOR_g NOR_1189_(.A(_0103_), .B(T2colour[2]), .Y(_0112_));
 NOR_g NOR_1190_(.A(_0112_), .B(_0111_), .Y(_0074_));
 NOR_g NOR_1253_(.A(T3state[0]), .B(T3state[1]), .Y(_0236_));
 NOR_g NOR_1260_(.A(T3y[1]), .B(T3y[0]), .Y(_0243_));
 NOR_g NOR_1263_(.A(_0244_), .B(T3y[3]), .Y(_0246_));
 NOR_g NOR_1267_(.A(_0248_), .B(T3y[6]), .Y(_0250_));
 NOR_g NOR_1272_(.A(_0254_), .B(_0250_), .Y(_0255_));
 NOR_g NOR_1273_(.A(_0255_), .B(_0242_), .Y(_0256_));
 NOR_g NOR_1274_(.A(T2Done), .B(T3state[3]), .Y(_0257_));
 NOR_g NOR_1275_(.A(_0257_), .B(_0256_), .Y(_0156_));
 NOR_g NOR_1277_(.A(T3state[2]), .B(T3state[3]), .Y(_0259_));
 NOR_g NOR_1284_(.A(_0265_), .B(_0262_), .Y(_0266_));
 NOR_g NOR_1317_(.A(_0296_), .B(T3x[7]), .Y(_0297_));
 NOR_g NOR_1323_(.A(T3plot), .B(KEY_N[0]), .Y(keywire1117));
 NOR_g NOR_1327_(.A(_0305_), .B(_0302_), .Y(_0306_));
 NOR_g NOR_1333_(.A(T3d[5]), .B(T3d[4]), .Y(_0311_));
 NOR_g NOR_1334_(.A(T3d[7]), .B(T3d[6]), .Y(_0312_));
 NOR_g NOR_1336_(.A(T3d[3]), .B(T3d[2]), .Y(_0314_));
 NOR_g NOR_1337_(.A(T3d[1]), .B(T3d[0]), .Y(_0315_));
 NOR_g NOR_1343_(.A(_0320_), .B(_0301_), .Y(_0321_));
 NOR_g NOR_1349_(.A(_0326_), .B(T3plot), .Y(_0327_));
 NOR_g NOR_1352_(.A(_0329_), .B(_0327_), .Y(_0330_));
 NOR_g NOR_1415_(.A(_0305_), .B(_0260_), .Y(_0383_));
 NOR_g NOR_1418_(.A(_0385_), .B(_0383_), .Y(_0386_));
 NOR_g NOR_1422_(.A(_0389_), .B(_0386_), .Y(_0390_));
 NOR_g NOR_1529_(.A(_0492_), .B(_0489_), .Y(_0493_));
 NOR_g NOR_1532_(.A(_0495_), .B(_0493_), .Y(_0496_));
 NOR_g NOR_1536_(.A(_0499_), .B(_0496_), .Y(_0500_));
 NOR_g NOR_1644_(.A(_0301_), .B(T3d[0]), .Y(_0604_));
 NOR_g NOR_1649_(.A(_0607_), .B(_0606_), .Y(_0608_));
 NOR_g NOR_1689_(.A(_0645_), .B(_0318_), .Y(_0646_));
 NOR_g NOR_1690_(.A(_0646_), .B(_0296_), .Y(_0647_));
 NOR_g NOR_1697_(.A(_0653_), .B(_0652_), .Y(_0654_));
 NOR_g NOR_1698_(.A(_0654_), .B(_0651_), .Y(_0655_));
 NOR_g NOR_1722_(.A(_0675_), .B(_0644_), .Y(_0678_));
 NOR_g NOR_1723_(.A(_0678_), .B(_0318_), .Y(_0679_));
 NOR_g NOR_1786_(.A(_0737_), .B(_0708_), .Y(_0740_));
 NOR_g NOR_1787_(.A(_0740_), .B(_0318_), .Y(_0741_));
 NOR_g NOR_1817_(.A(_0769_), .B(_0738_), .Y(_0770_));
 NOR_g NOR_1819_(.A(_0770_), .B(_0318_), .Y(_0772_));
 NOR_g NOR_1875_(.A(_0817_), .B(_0383_), .Y(_0818_));
 NOR_g NOR_1877_(.A(_0819_), .B(_0818_), .Y(_0820_));
 NOR_g NOR_1881_(.A(_0327_), .B(1'h1), .Y(_0824_));
 NOR_g NOR_1883_(.A(_0825_), .B(_0824_), .Y(_0826_));
 NOR_g NOR_1884_(.A(_0826_), .B(_0823_), .Y(_0827_));
 NOR_g NOR_1959_(.A(_0349_), .B(_0234_), .Y(_0899_));
 NOR_g NOR_1988_(.A(_0927_), .B(_0919_), .Y(_0928_));
 NOR_g NOR_1992_(.A(_0931_), .B(_0906_), .Y(_0932_));
 NOR_g NOR_1997_(.A(_0932_), .B(_0928_), .Y(_0937_));
 NOR_g NOR_2004_(.A(_0899_), .B(_0898_), .Y(_0943_));
 NOR_g NOR_2005_(.A(_0943_), .B(_0900_), .Y(_0944_));
 NOR_g NOR_2032_(.A(_0970_), .B(_0949_), .Y(_0971_));
 NOR_g NOR_2035_(.A(_0973_), .B(_0971_), .Y(_0974_));
 NOR_g NOR_2039_(.A(_0977_), .B(_0959_), .Y(_0978_));
 NOR_g NOR_2041_(.A(_0978_), .B(_0382_), .Y(_0980_));
 NOR_g NOR_2044_(.A(_0982_), .B(_0974_), .Y(_0983_));
 NOR_g NOR_2048_(.A(_0359_), .B(_0235_), .Y(_0986_));
 NOR_g NOR_2082_(.A(_1018_), .B(_0986_), .Y(_1019_));
 NOR_g NOR_2096_(.A(_1031_), .B(_1029_), .Y(_1033_));
 NOR_g NOR_2098_(.A(_1034_), .B(_1033_), .Y(_1035_));
 NOR_g NOR_2109_(.A(_0206_), .B(_1035_), .Y(_0207_));
 XOR_g XOR_1133_(.A(_0135_), .B(T2y[5]), .Y(_0146_));
 XOR_g XOR_1137_(.A(_0134_), .B(T2y[4]), .Y(_0075_));
 XOR_g XOR_1141_(.A(_0125_), .B(T2y[3]), .Y(_0078_));
 XOR_g XOR_1145_(.A(_0124_), .B(T2y[2]), .Y(_0081_));
 XOR_g XOR_1149_(.A(T2y[0]), .B(T2y[1]), .Y(_0084_));
 XOR_g XOR_1164_(.A(_0118_), .B(T2x[4]), .Y(keywire1168));
 XOR_g XOR_1167_(.A(_0117_), .B(T2x[3]), .Y(keywire1165));
 XOR_g XOR_1170_(.A(_0116_), .B(T2x[2]), .Y(keywire1162));
 XOR_g XOR_1173_(.A(T2x[0]), .B(T2x[1]), .Y(keywire1158));
 XOR_g XOR_1282_(.A(T3state[0]), .B(T3state[1]), .Y(_0264_));
 XOR_g XOR_1411_(.A(1'h1), .B(T3y[0]), .Y(_0379_));
 XOR_g XOR_1425_(.A(1'h1), .B(T3y[1]), .Y(_0392_));
 XOR_g XOR_1435_(.A(1'h1), .B(T3x[1]), .Y(_0402_));
 XOR_g XOR_1455_(.A(1'h1), .B(T3y[2]), .Y(_0421_));
 XOR_g XOR_1471_(.A(1'h1), .B(T3x[2]), .Y(_0437_));
 XOR_g XOR_1494_(.A(1'h1), .B(T3y[3]), .Y(_0459_));
 XOR_g XOR_1503_(.A(_0467_), .B(_0465_), .Y(_0468_));
 XOR_g XOR_1507_(.A(_0471_), .B(_0459_), .Y(_0472_));
 XOR_g XOR_1510_(.A(_0474_), .B(_0465_), .Y(_0475_));
 XOR_g XOR_1517_(.A(1'h0), .B(T3y[4]), .Y(_0481_));
 XOR_g XOR_1525_(.A(1'h0), .B(T3x[4]), .Y(_0489_));
 XOR_g XOR_1558_(.A(1'h0), .B(T3x[5]), .Y(_0521_));
 XOR_g XOR_1564_(.A(1'h0), .B(T3y[5]), .Y(_0527_));
 XOR_g XOR_1573_(.A(_0535_), .B(_0527_), .Y(_0536_));
 XOR_g XOR_1584_(.A(1'h1), .B(T3x[6]), .Y(_0546_));
 XOR_g XOR_1595_(.A(1'h1), .B(T3y[6]), .Y(_0557_));
 XOR_g XOR_1628_(.A(1'h0), .B(T3x[7]), .Y(_0589_));
 XOR_g XOR_1654_(.A(_0610_), .B(T3d[2]), .Y(_0612_));
 XOR_g XOR_1656_(.A(T3x[0]), .B(T3d[2]), .Y(_0614_));
 XOR_g XOR_1671_(.A(T3x[1]), .B(T3x[0]), .Y(_0628_));
 XOR_g XOR_1675_(.A(_0630_), .B(_0609_), .Y(_0632_));
 XOR_g XOR_1677_(.A(_0632_), .B(T3d[3]), .Y(_0634_));
 XOR_g XOR_1684_(.A(_0628_), .B(T3d[3]), .Y(_0641_));
 XOR_g XOR_1686_(.A(_0641_), .B(_0613_), .Y(_0643_));
 XOR_g XOR_1688_(.A(_0643_), .B(_0639_), .Y(_0645_));
 XOR_g XOR_1707_(.A(_0661_), .B(_0657_), .Y(_0663_));
 XOR_g XOR_1709_(.A(_0663_), .B(T3d[4]), .Y(_0665_));
 XOR_g XOR_1711_(.A(_0665_), .B(_0656_), .Y(_0667_));
 XOR_g XOR_1713_(.A(_0667_), .B(_0637_), .Y(_0669_));
 XOR_g XOR_1717_(.A(_0659_), .B(T3d[4]), .Y(_0673_));
 XOR_g XOR_1719_(.A(_0673_), .B(_0671_), .Y(_0675_));
 XOR_g XOR_1742_(.A(_0695_), .B(T3d[5]), .Y(_0697_));
 XOR_g XOR_1744_(.A(_0697_), .B(_0687_), .Y(_0699_));
 XOR_g XOR_1746_(.A(_0699_), .B(_0668_), .Y(_0701_));
 XOR_g XOR_1752_(.A(_0705_), .B(_0703_), .Y(_0707_));
 XOR_g XOR_1771_(.A(_0723_), .B(_0721_), .Y(_0725_));
 XOR_g XOR_1773_(.A(_0725_), .B(T3d[6]), .Y(_0727_));
 XOR_g XOR_1775_(.A(_0727_), .B(_0717_), .Y(_0729_));
 XOR_g XOR_1777_(.A(_0729_), .B(_0700_), .Y(_0731_));
 XOR_g XOR_1781_(.A(_0719_), .B(T3d[6]), .Y(_0735_));
 XOR_g XOR_1783_(.A(_0735_), .B(_0733_), .Y(_0737_));
 XOR_g XOR_1806_(.A(_0757_), .B(T3d[7]), .Y(_0759_));
 XOR_g XOR_1808_(.A(_0759_), .B(_0749_), .Y(_0761_));
 XOR_g XOR_1810_(.A(_0761_), .B(_0730_), .Y(_0763_));
 XOR_g XOR_1816_(.A(_0767_), .B(_0765_), .Y(_0769_));
 XOR_g XOR_1879_(.A(1'h1), .B(T3x[0]), .Y(_0822_));
 XOR_g XOR_1890_(.A(_0830_), .B(_0828_), .Y(_0832_));
 XOR_g XOR_1894_(.A(1'h1), .B(T3y[1]), .Y(_0836_));
 XOR_g XOR_1900_(.A(1'h1), .B(T3x[1]), .Y(_0842_));
 XOR_g XOR_1922_(.A(_0861_), .B(_0859_), .Y(_0863_));
 XOR_g XOR_1925_(.A(1'h0), .B(T3x[2]), .Y(_0866_));
 XOR_g XOR_1941_(.A(1'h0), .B(T3y[2]), .Y(_0882_));
 XOR_g XOR_1966_(.A(1'h1), .B(T3x[3]), .Y(_0906_));
 XOR_g XOR_1979_(.A(1'h1), .B(T3y[3]), .Y(_0919_));
 XOR_g XOR_2007_(.A(_0944_), .B(_0942_), .Y(_0946_));
 XOR_g XOR_2010_(.A(1'h1), .B(T3x[4]), .Y(_0949_));
 XOR_g XOR_2020_(.A(1'h1), .B(T3y[4]), .Y(_0959_));
 XOR_g XOR_2055_(.A(1'h1), .B(T3x[5]), .Y(_0993_));
 XOR_g XOR_2064_(.A(1'h1), .B(T3y[5]), .Y(_1002_));
 XOR_g XOR_2072_(.A(_1009_), .B(_0993_), .Y(_1010_));
 XOR_g XOR_2092_(.A(1'h0), .B(T3x[6]), .Y(_1029_));
 XOR_g keygate_XOR_2(.A(keywire1053), .B(lockingkeyinput[2]), .Y(T2x[1]));
 XOR_g keygate_XOR_3(.A(keywire1054), .B(lockingkeyinput[3]), .Y(T2x[2]));
 XOR_g keygate_XOR_4(.A(keywire1055), .B(lockingkeyinput[4]), .Y(T2x[3]));
 XOR_g keygate_XOR_7(.A(keywire1058), .B(lockingkeyinput[7]), .Y(T2x[6]));
 XOR_g keygate_XOR_8(.A(keywire1059), .B(lockingkeyinput[8]), .Y(T2x[7]));
 XOR_g keygate_XOR_15(.A(keywire1066), .B(lockingkeyinput[15]), .Y(T2y[6]));
 XOR_g keygate_XOR_17(.A(keywire1068), .B(lockingkeyinput[17]), .Y(T3state[0]));
 XOR_g keygate_XOR_18(.A(keywire1069), .B(lockingkeyinput[18]), .Y(T3state[1]));
 XOR_g keygate_XOR_19(.A(keywire1070), .B(lockingkeyinput[19]), .Y(T3state[2]));
 XOR_g keygate_XOR_20(.A(keywire1071), .B(lockingkeyinput[20]), .Y(T3state[3]));
 XOR_g keygate_XOR_24(.A(keywire1075), .B(lockingkeyinput[24]), .Y(T3y[0]));
 XOR_g keygate_XOR_25(.A(keywire1076), .B(lockingkeyinput[25]), .Y(T3y[1]));
 XOR_g keygate_XOR_26(.A(keywire1077), .B(lockingkeyinput[26]), .Y(T3y[2]));
 XOR_g keygate_XOR_28(.A(keywire1079), .B(lockingkeyinput[28]), .Y(T3y[4]));
 XOR_g keygate_XOR_30(.A(keywire1081), .B(lockingkeyinput[30]), .Y(T3y[6]));
 XOR_g keygate_XOR_31(.A(keywire1082), .B(lockingkeyinput[31]), .Y(T3colourcircle[0]));
 XOR_g keygate_XOR_34(.A(keywire1085), .B(lockingkeyinput[34]), .Y(T3xp[0]));
 XOR_g keygate_XOR_41(.A(keywire1092), .B(lockingkeyinput[41]), .Y(T3xp[7]));
 XOR_g keygate_XOR_42(.A(keywire1093), .B(lockingkeyinput[42]), .Y(T3d[0]));
 XOR_g keygate_XOR_46(.A(keywire1097), .B(lockingkeyinput[46]), .Y(T3d[4]));
 XOR_g keygate_XOR_48(.A(keywire1099), .B(lockingkeyinput[48]), .Y(T3d[6]));
 XOR_g keygate_XOR_49(.A(keywire1100), .B(lockingkeyinput[49]), .Y(T3d[7]));
 XOR_g keygate_XOR_50(.A(keywire1101), .B(lockingkeyinput[50]), .Y(T3d[8]));
 XOR_g keygate_XOR_52(.A(keywire1103), .B(lockingkeyinput[52]), .Y(T3x[1]));
 XOR_g keygate_XOR_53(.A(keywire1104), .B(lockingkeyinput[53]), .Y(T3x[2]));
 XOR_g keygate_XOR_55(.A(keywire1106), .B(lockingkeyinput[55]), .Y(T3x[4]));
 XOR_g keygate_XOR_56(.A(keywire1107), .B(lockingkeyinput[56]), .Y(T3x[5]));
 XOR_g keygate_XOR_57(.A(keywire1108), .B(lockingkeyinput[57]), .Y(T3x[6]));
 XOR_g keygate_XOR_58(.A(keywire1109), .B(lockingkeyinput[58]), .Y(T3x[7]));
 XOR_g keygate_XOR_63(.A(keywire1114), .B(lockingkeyinput[63]), .Y(T3yp[4]));
 XOR_g keygate_XOR_65(.A(keywire1116), .B(lockingkeyinput[65]), .Y(T3yp[6]));
 XOR_g keygate_XOR_71(.A(keywire1122), .B(lockingkeyinput[71]), .Y(_0044_));
 XOR_g keygate_XOR_72(.A(keywire1123), .B(lockingkeyinput[72]), .Y(_0045_));
 XOR_g keygate_XOR_73(.A(keywire1124), .B(lockingkeyinput[73]), .Y(_0046_));
 XOR_g keygate_XOR_75(.A(keywire1126), .B(lockingkeyinput[75]), .Y(_0048_));
 XOR_g keygate_XOR_77(.A(keywire1128), .B(lockingkeyinput[77]), .Y(_0050_));
 XOR_g keygate_XOR_78(.A(keywire1129), .B(lockingkeyinput[78]), .Y(_0051_));
 XOR_g keygate_XOR_79(.A(keywire1130), .B(lockingkeyinput[79]), .Y(_0052_));
 XOR_g keygate_XOR_81(.A(keywire1132), .B(lockingkeyinput[81]), .Y(_0054_));
 XOR_g keygate_XOR_82(.A(keywire1133), .B(lockingkeyinput[82]), .Y(_0055_));
 XOR_g keygate_XOR_83(.A(keywire1134), .B(lockingkeyinput[83]), .Y(_0149_));
 XOR_g keygate_XOR_84(.A(keywire1135), .B(lockingkeyinput[84]), .Y(_0150_));
 XOR_g keygate_XOR_86(.A(keywire1137), .B(lockingkeyinput[86]), .Y(_0152_));
 XOR_g keygate_XOR_88(.A(keywire1139), .B(lockingkeyinput[88]), .Y(_0368_));
 XOR_g keygate_XOR_89(.A(keywire1140), .B(lockingkeyinput[89]), .Y(_0370_));
 XOR_g keygate_XOR_91(.A(keywire1142), .B(lockingkeyinput[91]), .Y(_0228_));
 XOR_g keygate_XOR_92(.A(keywire1143), .B(lockingkeyinput[92]), .Y(_0229_));
 XOR_g keygate_XOR_93(.A(keywire1144), .B(lockingkeyinput[93]), .Y(_0653_));
 XOR_g keygate_XOR_94(.A(keywire1145), .B(lockingkeyinput[94]), .Y(_0323_));
 XOR_g keygate_XOR_95(.A(keywire1146), .B(lockingkeyinput[95]), .Y(_0341_));
 XOR_g keygate_XOR_97(.A(keywire1148), .B(lockingkeyinput[97]), .Y(_0356_));
 XOR_g keygate_XOR_98(.A(keywire1149), .B(lockingkeyinput[98]), .Y(_0324_));
 XOR_g keygate_XOR_100(.A(keywire1151), .B(lockingkeyinput[100]), .Y(_0359_));
 XOR_g keygate_XOR_107(.A(keywire1158), .B(lockingkeyinput[107]), .Y(_0100_));
 XOR_g keygate_XOR_108(.A(keywire1159), .B(lockingkeyinput[108]), .Y(_0037_));
 XOR_g keygate_XOR_112(.A(keywire1163), .B(lockingkeyinput[112]), .Y(_0002_));
 XOR_g keygate_XOR_113(.A(keywire1164), .B(lockingkeyinput[113]), .Y(_0118_));
 XOR_g keygate_XOR_114(.A(keywire1165), .B(lockingkeyinput[114]), .Y(_0096_));
 XOR_g keygate_XOR_120(.A(keywire1171), .B(lockingkeyinput[120]), .Y(_0120_));
 XOR_g keygate_XOR_122(.A(keywire1173), .B(lockingkeyinput[122]), .Y(_0115_));
 XOR_g keygate_XOR_124(.A(keywire1175), .B(lockingkeyinput[124]), .Y(_0090_));
 XOR_g keygate_XOR_126(.A(keywire1177), .B(lockingkeyinput[126]), .Y(_0114_));
 BUF_g BUF_1206_(.A(_0039_), .Y(T2Done));
 XNOR_g XNOR_1355_(.A(T3y[1]), .B(T3y[0]), .Y(_0332_));
 XNOR_g XNOR_1388_(.A(_0247_), .B(_0218_), .Y(_0361_));
 XNOR_g XNOR_1417_(.A(1'h1), .B(T3x[0]), .Y(_0385_));
 XNOR_g XNOR_1426_(.A(1'h1), .B(T3y[1]), .Y(_0393_));
 XNOR_g XNOR_1429_(.A(_0394_), .B(_0392_), .Y(_0396_));
 XNOR_g XNOR_1436_(.A(1'h1), .B(T3x[1]), .Y(_0403_));
 XNOR_g XNOR_1438_(.A(_0402_), .B(_0384_), .Y(_0405_));
 XNOR_g XNOR_1456_(.A(1'h1), .B(T3y[2]), .Y(_0422_));
 XNOR_g XNOR_1459_(.A(_0423_), .B(_0422_), .Y(_0425_));
 XNOR_g XNOR_1468_(.A(_0432_), .B(_0421_), .Y(_0434_));
 XNOR_g XNOR_1472_(.A(1'h1), .B(T3x[2]), .Y(_0438_));
 XNOR_g XNOR_1496_(.A(_0460_), .B(_0459_), .Y(_0461_));
 XNOR_g XNOR_1500_(.A(1'h1), .B(T3x[3]), .Y(_0465_));
 XNOR_g XNOR_1518_(.A(1'h0), .B(T3y[4]), .Y(_0482_));
 XNOR_g XNOR_1522_(.A(_0484_), .B(_0482_), .Y(_0486_));
 XNOR_g XNOR_1526_(.A(1'h0), .B(T3x[4]), .Y(_0490_));
 XNOR_g XNOR_1552_(.A(_0514_), .B(_0481_), .Y(_0516_));
 XNOR_g XNOR_1566_(.A(_0528_), .B(_0527_), .Y(_0529_));
 XNOR_g XNOR_1576_(.A(_0524_), .B(_0521_), .Y(_0539_));
 XNOR_g XNOR_1578_(.A(_0523_), .B(_0521_), .Y(_0541_));
 XNOR_g XNOR_1585_(.A(1'h1), .B(T3x[6]), .Y(_0547_));
 XNOR_g XNOR_1589_(.A(_0549_), .B(_0547_), .Y(_0551_));
 XNOR_g XNOR_1596_(.A(1'h1), .B(T3y[6]), .Y(_0558_));
 XNOR_g XNOR_1600_(.A(_0560_), .B(_0558_), .Y(_0562_));
 XNOR_g XNOR_1609_(.A(_0569_), .B(_0557_), .Y(_0571_));
 XNOR_g XNOR_1623_(.A(_0583_), .B(1'h0), .Y(_0584_));
 XNOR_g XNOR_1630_(.A(_0590_), .B(_0589_), .Y(_0591_));
 XNOR_g XNOR_1634_(.A(_0594_), .B(_0589_), .Y(_0595_));
 XNOR_g XNOR_1638_(.A(_0598_), .B(1'h0), .Y(_0599_));
 XNOR_g XNOR_1652_(.A(T3x[0]), .B(T3y[0]), .Y(_0610_));
 XNOR_g XNOR_1673_(.A(_0628_), .B(T3y[1]), .Y(_0630_));
 XNOR_g XNOR_1679_(.A(_0634_), .B(_0611_), .Y(_0636_));
 XNOR_g XNOR_1703_(.A(_0627_), .B(_0223_), .Y(_0659_));
 XNOR_g XNOR_1705_(.A(_0659_), .B(T3y[2]), .Y(_0661_));
 XNOR_g XNOR_1729_(.A(_0652_), .B(_0349_), .Y(_0685_));
 XNOR_g XNOR_1735_(.A(_0658_), .B(_0224_), .Y(_0690_));
 XNOR_g XNOR_1736_(.A(_0658_), .B(T3x[3]), .Y(_0691_));
 XNOR_g XNOR_1739_(.A(_0690_), .B(_0216_), .Y(_0694_));
 XNOR_g XNOR_1740_(.A(_0694_), .B(_0688_), .Y(_0695_));
 XNOR_g XNOR_1750_(.A(_0691_), .B(T3d[5]), .Y(_0705_));
 XNOR_g XNOR_1754_(.A(_0707_), .B(_0677_), .Y(_0709_));
 XNOR_g XNOR_1760_(.A(_0684_), .B(_0356_), .Y(_0715_));
 XNOR_g XNOR_1765_(.A(_0689_), .B(_0225_), .Y(_0719_));
 XNOR_g XNOR_1767_(.A(_0719_), .B(T3y[4]), .Y(_0721_));
 XNOR_g XNOR_1793_(.A(_0714_), .B(_0359_), .Y(_0747_));
 XNOR_g XNOR_1799_(.A(_0718_), .B(_0226_), .Y(_0752_));
 XNOR_g XNOR_1800_(.A(_0718_), .B(T3x[5]), .Y(_0753_));
 XNOR_g XNOR_1803_(.A(_0752_), .B(_0218_), .Y(_0756_));
 XNOR_g XNOR_1804_(.A(_0756_), .B(_0750_), .Y(_0757_));
 XNOR_g XNOR_1814_(.A(_0753_), .B(T3d[7]), .Y(_0767_));
 XNOR_g XNOR_1830_(.A(_0751_), .B(_0227_), .Y(_0782_));
 XNOR_g XNOR_1831_(.A(_0782_), .B(T3d[8]), .Y(_0783_));
 XNOR_g XNOR_1832_(.A(_0783_), .B(_0219_), .Y(_0784_));
 XNOR_g XNOR_1833_(.A(_0784_), .B(_0780_), .Y(_0785_));
 XNOR_g XNOR_1834_(.A(_0785_), .B(_0778_), .Y(_0786_));
 XNOR_g XNOR_1835_(.A(_0786_), .B(_0762_), .Y(_0787_));
 XNOR_g XNOR_1838_(.A(_0789_), .B(_0783_), .Y(_0790_));
 XNOR_g XNOR_1839_(.A(_0790_), .B(_0771_), .Y(_0791_));
 XNOR_g XNOR_1874_(.A(1'h1), .B(T3y[0]), .Y(_0817_));
 XNOR_g XNOR_1888_(.A(_0335_), .B(1'h1), .Y(_0830_));
 XNOR_g XNOR_1895_(.A(1'h1), .B(T3y[1]), .Y(_0837_));
 XNOR_g XNOR_1897_(.A(_0837_), .B(_0815_), .Y(_0839_));
 XNOR_g XNOR_1901_(.A(1'h1), .B(T3x[1]), .Y(_0843_));
 XNOR_g XNOR_1903_(.A(_0843_), .B(_0821_), .Y(_0845_));
 XNOR_g XNOR_1906_(.A(_0836_), .B(_0816_), .Y(_0848_));
 XNOR_g XNOR_1911_(.A(_0851_), .B(_0842_), .Y(_0853_));
 XNOR_g XNOR_1920_(.A(_0343_), .B(1'h0), .Y(_0861_));
 XNOR_g XNOR_1926_(.A(1'h0), .B(T3x[2]), .Y(_0867_));
 XNOR_g XNOR_1938_(.A(_0877_), .B(_0866_), .Y(_0879_));
 XNOR_g XNOR_1942_(.A(1'h0), .B(T3y[2]), .Y(_0883_));
 XNOR_g XNOR_1946_(.A(_0885_), .B(_0882_), .Y(_0887_));
 XNOR_g XNOR_1961_(.A(_0349_), .B(_0234_), .Y(_0901_));
 XNOR_g XNOR_1962_(.A(_0901_), .B(_0898_), .Y(_0902_));
 XNOR_g XNOR_2003_(.A(_0356_), .B(1'h1), .Y(_0942_));
 XNOR_g XNOR_2011_(.A(1'h1), .B(T3x[4]), .Y(_0950_));
 XNOR_g XNOR_2017_(.A(_0954_), .B(_0949_), .Y(_0956_));
 XNOR_g XNOR_2021_(.A(1'h1), .B(T3y[4]), .Y(_0960_));
 XNOR_g XNOR_2027_(.A(_0964_), .B(_0959_), .Y(_0966_));
 XNOR_g XNOR_2050_(.A(_0359_), .B(_0235_), .Y(_0988_));
 XNOR_g XNOR_2051_(.A(_0988_), .B(_0985_), .Y(_0989_));
 XNOR_g XNOR_2057_(.A(_0994_), .B(_0993_), .Y(_0995_));
 XNOR_g XNOR_2066_(.A(_1003_), .B(_1002_), .Y(_1004_));
 XNOR_g XNOR_2076_(.A(_1013_), .B(_1002_), .Y(_1014_));
 XNOR_g XNOR_2083_(.A(_1019_), .B(1'h0), .Y(_1020_));
 XNOR_g XNOR_2087_(.A(1'h0), .B(T3y[6]), .Y(_1024_));
 XNOR_g XNOR_2088_(.A(_1024_), .B(_1023_), .Y(_1025_));
 XNOR_g XNOR_2101_(.A(_1037_), .B(_1024_), .Y(_0199_));
 XNOR_g XNOR_2107_(.A(_0204_), .B(_1029_), .Y(_0205_));
 XNOR_g keygate_XNOR_0(.A(keywire1051), .B(lockingkeyinput[0]), .Y(vga_x[5]));
 XNOR_g keygate_XNOR_1(.A(keywire1052), .B(lockingkeyinput[1]), .Y(T2x[0]));
 XNOR_g keygate_XNOR_5(.A(keywire1056), .B(lockingkeyinput[5]), .Y(T2x[4]));
 XNOR_g keygate_XNOR_6(.A(keywire1057), .B(lockingkeyinput[6]), .Y(T2x[5]));
 XNOR_g keygate_XNOR_9(.A(keywire1060), .B(lockingkeyinput[9]), .Y(T2y[0]));
 XNOR_g keygate_XNOR_10(.A(keywire1061), .B(lockingkeyinput[10]), .Y(T2y[1]));
 XNOR_g keygate_XNOR_11(.A(keywire1062), .B(lockingkeyinput[11]), .Y(T2y[2]));
 XNOR_g keygate_XNOR_12(.A(keywire1063), .B(lockingkeyinput[12]), .Y(T2y[3]));
 XNOR_g keygate_XNOR_13(.A(keywire1064), .B(lockingkeyinput[13]), .Y(T2y[4]));
 XNOR_g keygate_XNOR_14(.A(keywire1065), .B(lockingkeyinput[14]), .Y(T2y[5]));
 XNOR_g keygate_XNOR_16(.A(keywire1067), .B(lockingkeyinput[16]), .Y(_0039_));
 XNOR_g keygate_XNOR_21(.A(keywire1072), .B(lockingkeyinput[21]), .Y(T2colour[0]));
 XNOR_g keygate_XNOR_22(.A(keywire1073), .B(lockingkeyinput[22]), .Y(T2colour[1]));
 XNOR_g keygate_XNOR_23(.A(keywire1074), .B(lockingkeyinput[23]), .Y(T2colour[2]));
 XNOR_g keygate_XNOR_27(.A(keywire1078), .B(lockingkeyinput[27]), .Y(T3y[3]));
 XNOR_g keygate_XNOR_29(.A(keywire1080), .B(lockingkeyinput[29]), .Y(T3y[5]));
 XNOR_g keygate_XNOR_32(.A(keywire1083), .B(lockingkeyinput[32]), .Y(T3colourcircle[1]));
 XNOR_g keygate_XNOR_33(.A(keywire1084), .B(lockingkeyinput[33]), .Y(T3colourcircle[2]));
 XNOR_g keygate_XNOR_35(.A(keywire1086), .B(lockingkeyinput[35]), .Y(T3xp[1]));
 XNOR_g keygate_XNOR_36(.A(keywire1087), .B(lockingkeyinput[36]), .Y(T3xp[2]));
 XNOR_g keygate_XNOR_37(.A(keywire1088), .B(lockingkeyinput[37]), .Y(T3xp[3]));
 XNOR_g keygate_XNOR_38(.A(keywire1089), .B(lockingkeyinput[38]), .Y(T3xp[4]));
 XNOR_g keygate_XNOR_39(.A(keywire1090), .B(lockingkeyinput[39]), .Y(T3xp[5]));
 XNOR_g keygate_XNOR_40(.A(keywire1091), .B(lockingkeyinput[40]), .Y(T3xp[6]));
 XNOR_g keygate_XNOR_43(.A(keywire1094), .B(lockingkeyinput[43]), .Y(T3d[1]));
 XNOR_g keygate_XNOR_44(.A(keywire1095), .B(lockingkeyinput[44]), .Y(T3d[2]));
 XNOR_g keygate_XNOR_45(.A(keywire1096), .B(lockingkeyinput[45]), .Y(T3d[3]));
 XNOR_g keygate_XNOR_47(.A(keywire1098), .B(lockingkeyinput[47]), .Y(T3d[5]));
 XNOR_g keygate_XNOR_51(.A(keywire1102), .B(lockingkeyinput[51]), .Y(T3x[0]));
 XNOR_g keygate_XNOR_54(.A(keywire1105), .B(lockingkeyinput[54]), .Y(T3x[3]));
 XNOR_g keygate_XNOR_59(.A(keywire1110), .B(lockingkeyinput[59]), .Y(T3yp[0]));
 XNOR_g keygate_XNOR_60(.A(keywire1111), .B(lockingkeyinput[60]), .Y(T3yp[1]));
 XNOR_g keygate_XNOR_61(.A(keywire1112), .B(lockingkeyinput[61]), .Y(T3yp[2]));
 XNOR_g keygate_XNOR_62(.A(keywire1113), .B(lockingkeyinput[62]), .Y(T3yp[3]));
 XNOR_g keygate_XNOR_64(.A(keywire1115), .B(lockingkeyinput[64]), .Y(T3yp[5]));
 XNOR_g keygate_XNOR_66(.A(keywire1117), .B(lockingkeyinput[66]), .Y(_0302_));
 XNOR_g keygate_XNOR_67(.A(keywire1118), .B(lockingkeyinput[67]), .Y(_0040_));
 XNOR_g keygate_XNOR_68(.A(keywire1119), .B(lockingkeyinput[68]), .Y(_0041_));
 XNOR_g keygate_XNOR_69(.A(keywire1120), .B(lockingkeyinput[69]), .Y(_0042_));
 XNOR_g keygate_XNOR_70(.A(keywire1121), .B(lockingkeyinput[70]), .Y(_0043_));
 XNOR_g keygate_XNOR_74(.A(keywire1125), .B(lockingkeyinput[74]), .Y(_0047_));
 XNOR_g keygate_XNOR_76(.A(keywire1127), .B(lockingkeyinput[76]), .Y(_0049_));
 XNOR_g keygate_XNOR_80(.A(keywire1131), .B(lockingkeyinput[80]), .Y(_0053_));
 XNOR_g keygate_XNOR_85(.A(keywire1136), .B(lockingkeyinput[85]), .Y(_0151_));
 XNOR_g keygate_XNOR_87(.A(keywire1138), .B(lockingkeyinput[87]), .Y(_0103_));
 XNOR_g keygate_XNOR_90(.A(keywire1141), .B(lockingkeyinput[90]), .Y(_0372_));
 XNOR_g keygate_XNOR_96(.A(keywire1147), .B(lockingkeyinput[96]), .Y(_0349_));
 XNOR_g keygate_XNOR_99(.A(keywire1150), .B(lockingkeyinput[99]), .Y(_0355_));
 XNOR_g keygate_XNOR_101(.A(keywire1152), .B(lockingkeyinput[101]), .Y(_0104_));
 XNOR_g keygate_XNOR_102(.A(keywire1153), .B(lockingkeyinput[102]), .Y(_0107_));
 XNOR_g keygate_XNOR_103(.A(keywire1154), .B(lockingkeyinput[103]), .Y(_0110_));
 XNOR_g keygate_XNOR_104(.A(keywire1155), .B(lockingkeyinput[104]), .Y(_0035_));
 XNOR_g keygate_XNOR_105(.A(keywire1156), .B(lockingkeyinput[105]), .Y(_0102_));
 XNOR_g keygate_XNOR_106(.A(keywire1157), .B(lockingkeyinput[106]), .Y(_0116_));
 XNOR_g keygate_XNOR_109(.A(keywire1160), .B(lockingkeyinput[109]), .Y(_0000_));
 XNOR_g keygate_XNOR_110(.A(keywire1161), .B(lockingkeyinput[110]), .Y(_0117_));
 XNOR_g keygate_XNOR_111(.A(keywire1162), .B(lockingkeyinput[111]), .Y(_0098_));
 XNOR_g keygate_XNOR_115(.A(keywire1166), .B(lockingkeyinput[115]), .Y(_0004_));
 XNOR_g keygate_XNOR_116(.A(keywire1167), .B(lockingkeyinput[116]), .Y(_0119_));
 XNOR_g keygate_XNOR_117(.A(keywire1168), .B(lockingkeyinput[117]), .Y(_0094_));
 XNOR_g keygate_XNOR_118(.A(keywire1169), .B(lockingkeyinput[118]), .Y(_0006_));
 XNOR_g keygate_XNOR_119(.A(keywire1170), .B(lockingkeyinput[119]), .Y(_0088_));
 XNOR_g keygate_XNOR_121(.A(keywire1172), .B(lockingkeyinput[121]), .Y(_0137_));
 XNOR_g keygate_XNOR_123(.A(keywire1174), .B(lockingkeyinput[123]), .Y(_0008_));
 XNOR_g keygate_XNOR_125(.A(keywire1176), .B(lockingkeyinput[125]), .Y(_0092_));
 XNOR_g keygate_XNOR_127(.A(keywire1178), .B(lockingkeyinput[127]), .Y(_0010_));
 DFFRcell DFF__1207_(.C(CLOCK_50), .D(_0056_), .Q(keywire1052), .R(_0040_));
 DFFRcell DFF__1208_(.C(CLOCK_50), .D(_0057_), .Q(keywire1053), .R(_0041_));
 DFFRcell DFF__1209_(.C(CLOCK_50), .D(_0058_), .Q(keywire1054), .R(_0042_));
 DFFRcell DFF__1210_(.C(CLOCK_50), .D(_0059_), .Q(keywire1055), .R(_0043_));
 DFFRcell DFF__1211_(.C(CLOCK_50), .D(_0060_), .Q(keywire1056), .R(_0044_));
 DFFRcell DFF__1212_(.C(CLOCK_50), .D(_0061_), .Q(keywire1057), .R(_0045_));
 DFFRcell DFF__1213_(.C(CLOCK_50), .D(_0062_), .Q(keywire1058), .R(_0046_));
 DFFRcell DFF__1214_(.C(CLOCK_50), .D(_0063_), .Q(keywire1059), .R(_0047_));
 DFFRcell DFF__1215_(.C(CLOCK_50), .D(_0064_), .Q(keywire1060), .R(_0048_));
 DFFRcell DFF__1216_(.C(CLOCK_50), .D(_0065_), .Q(keywire1061), .R(_0049_));
 DFFRcell DFF__1217_(.C(CLOCK_50), .D(_0066_), .Q(keywire1062), .R(_0050_));
 DFFRcell DFF__1218_(.C(CLOCK_50), .D(_0067_), .Q(keywire1063), .R(_0051_));
 DFFRcell DFF__1219_(.C(CLOCK_50), .D(_0068_), .Q(keywire1064), .R(_0052_));
 DFFRcell DFF__1220_(.C(CLOCK_50), .D(_0069_), .Q(keywire1065), .R(_0053_));
 DFFRcell DFF__1221_(.C(CLOCK_50), .D(_0070_), .Q(keywire1066), .R(_0054_));
 DFFRcell DFF__1222_(.C(CLOCK_50), .D(_0071_), .Q(keywire1067), .R(_0055_));
 DFFRcell DFF__2116_(.C(CLOCK_50), .D(_0153_), .Q(keywire1068), .R(_0149_));
 DFFRcell DFF__2117_(.C(CLOCK_50), .D(_0154_), .Q(keywire1069), .R(_0150_));
 DFFRcell DFF__2118_(.C(CLOCK_50), .D(_0155_), .Q(keywire1070), .R(_0151_));
 DFFRcell DFF__2119_(.C(CLOCK_50), .D(_0156_), .Q(keywire1071), .R(_0152_));
 DFFcell DFF__1223_(.C(CLOCK_50), .D(_0072_), .Q(keywire1072));
 DFFcell DFF__1224_(.C(CLOCK_50), .D(_0073_), .Q(keywire1073));
 DFFcell DFF__1225_(.C(CLOCK_50), .D(_0074_), .Q(keywire1074));
 DFFcell DFF__2120_(.C(CLOCK_50), .D(_0157_), .Q(keywire1075));
 DFFcell DFF__2121_(.C(CLOCK_50), .D(_0158_), .Q(keywire1076));
 DFFcell DFF__2122_(.C(CLOCK_50), .D(_0159_), .Q(keywire1077));
 DFFcell DFF__2123_(.C(CLOCK_50), .D(_0160_), .Q(keywire1078));
 DFFcell DFF__2124_(.C(CLOCK_50), .D(_0161_), .Q(keywire1079));
 DFFcell DFF__2125_(.C(CLOCK_50), .D(_0162_), .Q(keywire1080));
 DFFcell DFF__2126_(.C(CLOCK_50), .D(_0163_), .Q(keywire1081));
 DFFcell DFF__2127_(.C(CLOCK_50), .D(_0164_), .Q(keywire1082));
 DFFcell DFF__2128_(.C(CLOCK_50), .D(_0165_), .Q(keywire1083));
 DFFcell DFF__2129_(.C(CLOCK_50), .D(_0166_), .Q(keywire1084));
 DFFcell DFF__2130_(.C(CLOCK_50), .D(_0167_), .Q(keywire1085));
 DFFcell DFF__2131_(.C(CLOCK_50), .D(_0168_), .Q(keywire1086));
 DFFcell DFF__2132_(.C(CLOCK_50), .D(_0169_), .Q(keywire1087));
 DFFcell DFF__2133_(.C(CLOCK_50), .D(_0170_), .Q(keywire1088));
 DFFcell DFF__2134_(.C(CLOCK_50), .D(_0171_), .Q(keywire1089));
 DFFcell DFF__2135_(.C(CLOCK_50), .D(_0172_), .Q(keywire1090));
 DFFcell DFF__2136_(.C(CLOCK_50), .D(_0173_), .Q(keywire1091));
 DFFcell DFF__2137_(.C(CLOCK_50), .D(_0174_), .Q(keywire1092));
 DFFcell DFF__2138_(.C(CLOCK_50), .D(_0175_), .Q(keywire1093));
 DFFcell DFF__2139_(.C(CLOCK_50), .D(_0176_), .Q(keywire1094));
 DFFcell DFF__2140_(.C(CLOCK_50), .D(_0177_), .Q(keywire1095));
 DFFcell DFF__2141_(.C(CLOCK_50), .D(_0178_), .Q(keywire1096));
 DFFcell DFF__2142_(.C(CLOCK_50), .D(_0179_), .Q(keywire1097));
 DFFcell DFF__2143_(.C(CLOCK_50), .D(_0180_), .Q(keywire1098));
 DFFcell DFF__2144_(.C(CLOCK_50), .D(_0181_), .Q(keywire1099));
 DFFcell DFF__2145_(.C(CLOCK_50), .D(_0182_), .Q(keywire1100));
 DFFcell DFF__2146_(.C(CLOCK_50), .D(_0183_), .Q(keywire1101));
 DFFcell DFF__2147_(.C(CLOCK_50), .D(_0184_), .Q(keywire1102));
 DFFcell DFF__2148_(.C(CLOCK_50), .D(_0185_), .Q(keywire1103));
 DFFcell DFF__2149_(.C(CLOCK_50), .D(_0186_), .Q(keywire1104));
 DFFcell DFF__2150_(.C(CLOCK_50), .D(_0187_), .Q(keywire1105));
 DFFcell DFF__2151_(.C(CLOCK_50), .D(_0188_), .Q(keywire1106));
 DFFcell DFF__2152_(.C(CLOCK_50), .D(_0189_), .Q(keywire1107));
 DFFcell DFF__2153_(.C(CLOCK_50), .D(_0190_), .Q(keywire1108));
 DFFcell DFF__2154_(.C(CLOCK_50), .D(_0191_), .Q(keywire1109));
 DFFcell DFF__2155_(.C(CLOCK_50), .D(_0192_), .Q(keywire1110));
 DFFcell DFF__2156_(.C(CLOCK_50), .D(_0193_), .Q(keywire1111));
 DFFcell DFF__2157_(.C(CLOCK_50), .D(_0194_), .Q(keywire1112));
 DFFcell DFF__2158_(.C(CLOCK_50), .D(_0195_), .Q(keywire1113));
 DFFcell DFF__2159_(.C(CLOCK_50), .D(_0196_), .Q(keywire1114));
 DFFcell DFF__2160_(.C(CLOCK_50), .D(_0197_), .Q(keywire1115));
 DFFcell DFF__2161_(.C(CLOCK_50), .D(_0198_), .Q(keywire1116));
endmodule
 


module BUF_g(A, Y);
input A;
output Y;
assign Y=A;
endmodule

 
module NOT_g(A, Y);
input A;
output Y;
assign Y=~A;
endmodule

module AND_g(A, B, Y);
input A, B;
output Y;
assign Y=(A & B);
endmodule

module OR_g(A, B, Y);
input A, B;
output Y;
assign Y= (A | B);
endmodule

module NAND_g(A, B, Y);
input A, B;
output Y;
assign Y= ~(A & B);

endmodule

module NOR_g(A, B, Y);
input A, B;
output Y;
assign Y = ~(A | B);
endmodule


module XOR_g(A, B, Y);
input A, B;
output Y;
assign Y = (A ^ B);
endmodule

module XNOR_g(A, B, Y);
input A, B;
output Y;
assign Y = ~(A ^ B);
endmodule

module DFFcell(C, D, Q);
input C, D;
output reg Q;
always @(posedge C)
	Q <= D;
endmodule


module DFFRcell(C, D, Q, R);
input C, D, R;
wire x;
assign x=~R;
output reg Q;
always @(posedge C, negedge x)
	if (!x)
		Q <= 1'b0;
	else
		Q <= D;
endmodule
